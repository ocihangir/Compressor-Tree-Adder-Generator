// (* RLOC_ORIGIN = "X0Y0" *)
module mult_64x64_lut6(in0, in1, mult_out);

input [63:0] in0;
input [63:0] in1;
output [128:0] mult_out;

wire [63:0] pp0;
assign pp0 = (in1[0]) ? in0 : 1'b0;
wire [63:0] pp1;
assign pp1 = (in1[1]) ? in0 : 1'b0;
wire [63:0] pp2;
assign pp2 = (in1[2]) ? in0 : 1'b0;
wire [63:0] pp3;
assign pp3 = (in1[3]) ? in0 : 1'b0;
wire [63:0] pp4;
assign pp4 = (in1[4]) ? in0 : 1'b0;
wire [63:0] pp5;
assign pp5 = (in1[5]) ? in0 : 1'b0;
wire [63:0] pp6;
assign pp6 = (in1[6]) ? in0 : 1'b0;
wire [63:0] pp7;
assign pp7 = (in1[7]) ? in0 : 1'b0;
wire [63:0] pp8;
assign pp8 = (in1[8]) ? in0 : 1'b0;
wire [63:0] pp9;
assign pp9 = (in1[9]) ? in0 : 1'b0;
wire [63:0] pp10;
assign pp10 = (in1[10]) ? in0 : 1'b0;
wire [63:0] pp11;
assign pp11 = (in1[11]) ? in0 : 1'b0;
wire [63:0] pp12;
assign pp12 = (in1[12]) ? in0 : 1'b0;
wire [63:0] pp13;
assign pp13 = (in1[13]) ? in0 : 1'b0;
wire [63:0] pp14;
assign pp14 = (in1[14]) ? in0 : 1'b0;
wire [63:0] pp15;
assign pp15 = (in1[15]) ? in0 : 1'b0;
wire [63:0] pp16;
assign pp16 = (in1[16]) ? in0 : 1'b0;
wire [63:0] pp17;
assign pp17 = (in1[17]) ? in0 : 1'b0;
wire [63:0] pp18;
assign pp18 = (in1[18]) ? in0 : 1'b0;
wire [63:0] pp19;
assign pp19 = (in1[19]) ? in0 : 1'b0;
wire [63:0] pp20;
assign pp20 = (in1[20]) ? in0 : 1'b0;
wire [63:0] pp21;
assign pp21 = (in1[21]) ? in0 : 1'b0;
wire [63:0] pp22;
assign pp22 = (in1[22]) ? in0 : 1'b0;
wire [63:0] pp23;
assign pp23 = (in1[23]) ? in0 : 1'b0;
wire [63:0] pp24;
assign pp24 = (in1[24]) ? in0 : 1'b0;
wire [63:0] pp25;
assign pp25 = (in1[25]) ? in0 : 1'b0;
wire [63:0] pp26;
assign pp26 = (in1[26]) ? in0 : 1'b0;
wire [63:0] pp27;
assign pp27 = (in1[27]) ? in0 : 1'b0;
wire [63:0] pp28;
assign pp28 = (in1[28]) ? in0 : 1'b0;
wire [63:0] pp29;
assign pp29 = (in1[29]) ? in0 : 1'b0;
wire [63:0] pp30;
assign pp30 = (in1[30]) ? in0 : 1'b0;
wire [63:0] pp31;
assign pp31 = (in1[31]) ? in0 : 1'b0;
wire [63:0] pp32;
assign pp32 = (in1[32]) ? in0 : 1'b0;
wire [63:0] pp33;
assign pp33 = (in1[33]) ? in0 : 1'b0;
wire [63:0] pp34;
assign pp34 = (in1[34]) ? in0 : 1'b0;
wire [63:0] pp35;
assign pp35 = (in1[35]) ? in0 : 1'b0;
wire [63:0] pp36;
assign pp36 = (in1[36]) ? in0 : 1'b0;
wire [63:0] pp37;
assign pp37 = (in1[37]) ? in0 : 1'b0;
wire [63:0] pp38;
assign pp38 = (in1[38]) ? in0 : 1'b0;
wire [63:0] pp39;
assign pp39 = (in1[39]) ? in0 : 1'b0;
wire [63:0] pp40;
assign pp40 = (in1[40]) ? in0 : 1'b0;
wire [63:0] pp41;
assign pp41 = (in1[41]) ? in0 : 1'b0;
wire [63:0] pp42;
assign pp42 = (in1[42]) ? in0 : 1'b0;
wire [63:0] pp43;
assign pp43 = (in1[43]) ? in0 : 1'b0;
wire [63:0] pp44;
assign pp44 = (in1[44]) ? in0 : 1'b0;
wire [63:0] pp45;
assign pp45 = (in1[45]) ? in0 : 1'b0;
wire [63:0] pp46;
assign pp46 = (in1[46]) ? in0 : 1'b0;
wire [63:0] pp47;
assign pp47 = (in1[47]) ? in0 : 1'b0;
wire [63:0] pp48;
assign pp48 = (in1[48]) ? in0 : 1'b0;
wire [63:0] pp49;
assign pp49 = (in1[49]) ? in0 : 1'b0;
wire [63:0] pp50;
assign pp50 = (in1[50]) ? in0 : 1'b0;
wire [63:0] pp51;
assign pp51 = (in1[51]) ? in0 : 1'b0;
wire [63:0] pp52;
assign pp52 = (in1[52]) ? in0 : 1'b0;
wire [63:0] pp53;
assign pp53 = (in1[53]) ? in0 : 1'b0;
wire [63:0] pp54;
assign pp54 = (in1[54]) ? in0 : 1'b0;
wire [63:0] pp55;
assign pp55 = (in1[55]) ? in0 : 1'b0;
wire [63:0] pp56;
assign pp56 = (in1[56]) ? in0 : 1'b0;
wire [63:0] pp57;
assign pp57 = (in1[57]) ? in0 : 1'b0;
wire [63:0] pp58;
assign pp58 = (in1[58]) ? in0 : 1'b0;
wire [63:0] pp59;
assign pp59 = (in1[59]) ? in0 : 1'b0;
wire [63:0] pp60;
assign pp60 = (in1[60]) ? in0 : 1'b0;
wire [63:0] pp61;
assign pp61 = (in1[61]) ? in0 : 1'b0;
wire [63:0] pp62;
assign pp62 = (in1[62]) ? in0 : 1'b0;
wire [63:0] pp63;
assign pp63 = (in1[63]) ? in0 : 1'b0;
wire [2:0] gpcOutL1_0;

// (* RLOC = "X1Y0" *)
gpc006 gpcL1_0 ({pp0[63],pp1[62],pp2[61],pp3[60],pp4[59],pp5[58]},gpcOutL1_0);
wire [2:0] gpcOutL1_1;

// (* RLOC = "X1Y1" *)
gpc006 gpcL1_1 ({pp0[62],pp1[61],pp2[60],pp3[59],pp4[58],pp5[57]},gpcOutL1_1);
wire [2:0] gpcOutL1_2;

// (* RLOC = "X1Y2" *)
gpc006 gpcL1_2 ({pp1[63],pp2[62],pp3[61],pp4[60],pp5[59],pp6[58]},gpcOutL1_2);
wire [2:0] gpcOutL1_3;

// (* RLOC = "X1Y3" *)
gpc006 gpcL1_3 ({pp0[61],pp1[60],pp2[59],pp3[58],pp4[57],pp5[56]},gpcOutL1_3);
wire [2:0] gpcOutL1_4;

// (* RLOC = "X1Y4" *)
gpc006 gpcL1_4 ({pp2[63],pp3[62],pp4[61],pp5[60],pp6[59],pp7[58]},gpcOutL1_4);
wire [2:0] gpcOutL1_5;

// (* RLOC = "X1Y5" *)
gpc006 gpcL1_5 ({pp0[60],pp1[59],pp2[58],pp3[57],pp4[56],pp5[55]},gpcOutL1_5);
wire [2:0] gpcOutL1_6;

// (* RLOC = "X1Y6" *)
gpc006 gpcL1_6 ({pp3[63],pp4[62],pp5[61],pp6[60],pp7[59],pp8[58]},gpcOutL1_6);
wire [2:0] gpcOutL1_7;

// (* RLOC = "X1Y7" *)
gpc006 gpcL1_7 ({pp0[59],pp1[58],pp2[57],pp3[56],pp4[55],pp5[54]},gpcOutL1_7);
wire [2:0] gpcOutL1_8;

// (* RLOC = "X1Y8" *)
gpc006 gpcL1_8 ({pp4[63],pp5[62],pp6[61],pp7[60],pp8[59],pp9[58]},gpcOutL1_8);
wire [2:0] gpcOutL1_9;

// (* RLOC = "X1Y9" *)
gpc006 gpcL1_9 ({pp0[58],pp1[57],pp2[56],pp3[55],pp4[54],pp5[53]},gpcOutL1_9);
wire [2:0] gpcOutL1_10;

// (* RLOC = "X1Y10" *)
gpc006 gpcL1_10 ({pp5[63],pp6[62],pp7[61],pp8[60],pp9[59],pp10[58]},gpcOutL1_10);
wire [2:0] gpcOutL1_11;

// (* RLOC = "X1Y11" *)
gpc006 gpcL1_11 ({pp0[57],pp1[56],pp2[55],pp3[54],pp4[53],pp5[52]},gpcOutL1_11);
wire [2:0] gpcOutL1_12;

// (* RLOC = "X1Y12" *)
gpc006 gpcL1_12 ({pp6[57],pp7[56],pp8[55],pp9[54],pp10[53],pp11[52]},gpcOutL1_12);
wire [2:0] gpcOutL1_13;

// (* RLOC = "X1Y13" *)
gpc006 gpcL1_13 ({pp6[63],pp7[62],pp8[61],pp9[60],pp10[59],pp11[58]},gpcOutL1_13);
wire [2:0] gpcOutL1_14;

// (* RLOC = "X1Y14" *)
gpc006 gpcL1_14 ({pp0[56],pp1[55],pp2[54],pp3[53],pp4[52],pp5[51]},gpcOutL1_14);
wire [2:0] gpcOutL1_15;

// (* RLOC = "X1Y15" *)
gpc006 gpcL1_15 ({pp6[56],pp7[55],pp8[54],pp9[53],pp10[52],pp11[51]},gpcOutL1_15);
wire [2:0] gpcOutL1_16;

// (* RLOC = "X1Y16" *)
gpc006 gpcL1_16 ({pp7[57],pp8[56],pp9[55],pp10[54],pp11[53],pp12[52]},gpcOutL1_16);
wire [2:0] gpcOutL1_17;

// (* RLOC = "X1Y17" *)
gpc006 gpcL1_17 ({pp7[63],pp8[62],pp9[61],pp10[60],pp11[59],pp12[58]},gpcOutL1_17);
wire [2:0] gpcOutL1_18;

// (* RLOC = "X1Y18" *)
gpc006 gpcL1_18 ({pp0[55],pp1[54],pp2[53],pp3[52],pp4[51],pp5[50]},gpcOutL1_18);
wire [2:0] gpcOutL1_19;

// (* RLOC = "X1Y19" *)
gpc006 gpcL1_19 ({pp6[55],pp7[54],pp8[53],pp9[52],pp10[51],pp11[50]},gpcOutL1_19);
wire [2:0] gpcOutL1_20;

// (* RLOC = "X1Y20" *)
gpc006 gpcL1_20 ({pp8[57],pp9[56],pp10[55],pp11[54],pp12[53],pp13[52]},gpcOutL1_20);
wire [2:0] gpcOutL1_21;

// (* RLOC = "X1Y21" *)
gpc006 gpcL1_21 ({pp8[63],pp9[62],pp10[61],pp11[60],pp12[59],pp13[58]},gpcOutL1_21);
wire [2:0] gpcOutL1_22;

// (* RLOC = "X1Y22" *)
gpc006 gpcL1_22 ({pp0[54],pp1[53],pp2[52],pp3[51],pp4[50],pp5[49]},gpcOutL1_22);
wire [2:0] gpcOutL1_23;

// (* RLOC = "X1Y23" *)
gpc006 gpcL1_23 ({pp6[54],pp7[53],pp8[52],pp9[51],pp10[50],pp11[49]},gpcOutL1_23);
wire [2:0] gpcOutL1_24;

// (* RLOC = "X1Y24" *)
gpc006 gpcL1_24 ({pp9[57],pp10[56],pp11[55],pp12[54],pp13[53],pp14[52]},gpcOutL1_24);
wire [2:0] gpcOutL1_25;

// (* RLOC = "X1Y25" *)
gpc006 gpcL1_25 ({pp9[63],pp10[62],pp11[61],pp12[60],pp13[59],pp14[58]},gpcOutL1_25);
wire [2:0] gpcOutL1_26;

// (* RLOC = "X1Y26" *)
gpc006 gpcL1_26 ({pp0[53],pp1[52],pp2[51],pp3[50],pp4[49],pp5[48]},gpcOutL1_26);
wire [2:0] gpcOutL1_27;

// (* RLOC = "X1Y27" *)
gpc006 gpcL1_27 ({pp6[53],pp7[52],pp8[51],pp9[50],pp10[49],pp11[48]},gpcOutL1_27);
wire [2:0] gpcOutL1_28;

// (* RLOC = "X1Y28" *)
gpc006 gpcL1_28 ({pp10[57],pp11[56],pp12[55],pp13[54],pp14[53],pp15[52]},gpcOutL1_28);
wire [2:0] gpcOutL1_29;

// (* RLOC = "X1Y29" *)
gpc006 gpcL1_29 ({pp10[63],pp11[62],pp12[61],pp13[60],pp14[59],pp15[58]},gpcOutL1_29);
wire [2:0] gpcOutL1_30;

// (* RLOC = "X1Y30" *)
gpc006 gpcL1_30 ({pp0[52],pp1[51],pp2[50],pp3[49],pp4[48],pp5[47]},gpcOutL1_30);
wire [2:0] gpcOutL1_31;

// (* RLOC = "X1Y31" *)
gpc006 gpcL1_31 ({pp6[52],pp7[51],pp8[50],pp9[49],pp10[48],pp11[47]},gpcOutL1_31);
wire [2:0] gpcOutL1_32;

// (* RLOC = "X1Y32" *)
gpc006 gpcL1_32 ({pp11[57],pp12[56],pp13[55],pp14[54],pp15[53],pp16[52]},gpcOutL1_32);
wire [2:0] gpcOutL1_33;

// (* RLOC = "X1Y33" *)
gpc006 gpcL1_33 ({pp11[63],pp12[62],pp13[61],pp14[60],pp15[59],pp16[58]},gpcOutL1_33);
wire [2:0] gpcOutL1_34;

// (* RLOC = "X1Y34" *)
gpc006 gpcL1_34 ({pp0[51],pp1[50],pp2[49],pp3[48],pp4[47],pp5[46]},gpcOutL1_34);
wire [2:0] gpcOutL1_35;

// (* RLOC = "X1Y35" *)
gpc006 gpcL1_35 ({pp6[51],pp7[50],pp8[49],pp9[48],pp10[47],pp11[46]},gpcOutL1_35);
wire [2:0] gpcOutL1_36;

// (* RLOC = "X1Y36" *)
gpc006 gpcL1_36 ({pp12[51],pp13[50],pp14[49],pp15[48],pp16[47],pp17[46]},gpcOutL1_36);
wire [2:0] gpcOutL1_37;

// (* RLOC = "X1Y37" *)
gpc006 gpcL1_37 ({pp12[57],pp13[56],pp14[55],pp15[54],pp16[53],pp17[52]},gpcOutL1_37);
wire [2:0] gpcOutL1_38;

// (* RLOC = "X1Y38" *)
gpc006 gpcL1_38 ({pp12[63],pp13[62],pp14[61],pp15[60],pp16[59],pp17[58]},gpcOutL1_38);
wire [2:0] gpcOutL1_39;

// (* RLOC = "X1Y39" *)
gpc006 gpcL1_39 ({pp0[50],pp1[49],pp2[48],pp3[47],pp4[46],pp5[45]},gpcOutL1_39);
wire [2:0] gpcOutL1_40;

// (* RLOC = "X1Y40" *)
gpc006 gpcL1_40 ({pp6[50],pp7[49],pp8[48],pp9[47],pp10[46],pp11[45]},gpcOutL1_40);
wire [2:0] gpcOutL1_41;

// (* RLOC = "X1Y41" *)
gpc006 gpcL1_41 ({pp12[50],pp13[49],pp14[48],pp15[47],pp16[46],pp17[45]},gpcOutL1_41);
wire [2:0] gpcOutL1_42;

// (* RLOC = "X1Y42" *)
gpc006 gpcL1_42 ({pp13[51],pp14[50],pp15[49],pp16[48],pp17[47],pp18[46]},gpcOutL1_42);
wire [2:0] gpcOutL1_43;

// (* RLOC = "X1Y43" *)
gpc006 gpcL1_43 ({pp13[57],pp14[56],pp15[55],pp16[54],pp17[53],pp18[52]},gpcOutL1_43);
wire [2:0] gpcOutL1_44;

// (* RLOC = "X1Y44" *)
gpc006 gpcL1_44 ({pp13[63],pp14[62],pp15[61],pp16[60],pp17[59],pp18[58]},gpcOutL1_44);
wire [2:0] gpcOutL1_45;

// (* RLOC = "X1Y45" *)
gpc006 gpcL1_45 ({pp0[49],pp1[48],pp2[47],pp3[46],pp4[45],pp5[44]},gpcOutL1_45);
wire [2:0] gpcOutL1_46;

// (* RLOC = "X1Y46" *)
gpc006 gpcL1_46 ({pp6[49],pp7[48],pp8[47],pp9[46],pp10[45],pp11[44]},gpcOutL1_46);
wire [2:0] gpcOutL1_47;

// (* RLOC = "X1Y47" *)
gpc006 gpcL1_47 ({pp12[49],pp13[48],pp14[47],pp15[46],pp16[45],pp17[44]},gpcOutL1_47);
wire [2:0] gpcOutL1_48;

// (* RLOC = "X1Y48" *)
gpc006 gpcL1_48 ({pp14[51],pp15[50],pp16[49],pp17[48],pp18[47],pp19[46]},gpcOutL1_48);
wire [2:0] gpcOutL1_49;

// (* RLOC = "X1Y49" *)
gpc006 gpcL1_49 ({pp14[57],pp15[56],pp16[55],pp17[54],pp18[53],pp19[52]},gpcOutL1_49);
wire [2:0] gpcOutL1_50;

// (* RLOC = "X1Y50" *)
gpc006 gpcL1_50 ({pp14[63],pp15[62],pp16[61],pp17[60],pp18[59],pp19[58]},gpcOutL1_50);
wire [2:0] gpcOutL1_51;

// (* RLOC = "X1Y51" *)
gpc006 gpcL1_51 ({pp0[48],pp1[47],pp2[46],pp3[45],pp4[44],pp5[43]},gpcOutL1_51);
wire [2:0] gpcOutL1_52;

// (* RLOC = "X1Y52" *)
gpc006 gpcL1_52 ({pp6[48],pp7[47],pp8[46],pp9[45],pp10[44],pp11[43]},gpcOutL1_52);
wire [2:0] gpcOutL1_53;

// (* RLOC = "X1Y53" *)
gpc006 gpcL1_53 ({pp12[48],pp13[47],pp14[46],pp15[45],pp16[44],pp17[43]},gpcOutL1_53);
wire [2:0] gpcOutL1_54;

// (* RLOC = "X1Y54" *)
gpc006 gpcL1_54 ({pp15[51],pp16[50],pp17[49],pp18[48],pp19[47],pp20[46]},gpcOutL1_54);
wire [2:0] gpcOutL1_55;

// (* RLOC = "X1Y55" *)
gpc006 gpcL1_55 ({pp15[57],pp16[56],pp17[55],pp18[54],pp19[53],pp20[52]},gpcOutL1_55);
wire [2:0] gpcOutL1_56;

// (* RLOC = "X1Y56" *)
gpc006 gpcL1_56 ({pp15[63],pp16[62],pp17[61],pp18[60],pp19[59],pp20[58]},gpcOutL1_56);
wire [2:0] gpcOutL1_57;

// (* RLOC = "X1Y57" *)
gpc006 gpcL1_57 ({pp0[47],pp1[46],pp2[45],pp3[44],pp4[43],pp5[42]},gpcOutL1_57);
wire [2:0] gpcOutL1_58;

// (* RLOC = "X1Y58" *)
gpc006 gpcL1_58 ({pp6[47],pp7[46],pp8[45],pp9[44],pp10[43],pp11[42]},gpcOutL1_58);
wire [2:0] gpcOutL1_59;

// (* RLOC = "X1Y59" *)
gpc006 gpcL1_59 ({pp12[47],pp13[46],pp14[45],pp15[44],pp16[43],pp17[42]},gpcOutL1_59);
wire [2:0] gpcOutL1_60;

// (* RLOC = "X1Y60" *)
gpc006 gpcL1_60 ({pp16[51],pp17[50],pp18[49],pp19[48],pp20[47],pp21[46]},gpcOutL1_60);
wire [2:0] gpcOutL1_61;

// (* RLOC = "X1Y61" *)
gpc006 gpcL1_61 ({pp16[57],pp17[56],pp18[55],pp19[54],pp20[53],pp21[52]},gpcOutL1_61);
wire [2:0] gpcOutL1_62;

// (* RLOC = "X1Y62" *)
gpc006 gpcL1_62 ({pp16[63],pp17[62],pp18[61],pp19[60],pp20[59],pp21[58]},gpcOutL1_62);
wire [2:0] gpcOutL1_63;

// (* RLOC = "X1Y63" *)
gpc006 gpcL1_63 ({pp0[46],pp1[45],pp2[44],pp3[43],pp4[42],pp5[41]},gpcOutL1_63);
wire [2:0] gpcOutL1_64;

// (* RLOC = "X1Y64" *)
gpc006 gpcL1_64 ({pp6[46],pp7[45],pp8[44],pp9[43],pp10[42],pp11[41]},gpcOutL1_64);
wire [2:0] gpcOutL1_65;

// (* RLOC = "X1Y65" *)
gpc006 gpcL1_65 ({pp12[46],pp13[45],pp14[44],pp15[43],pp16[42],pp17[41]},gpcOutL1_65);
wire [2:0] gpcOutL1_66;

// (* RLOC = "X1Y66" *)
gpc006 gpcL1_66 ({pp17[51],pp18[50],pp19[49],pp20[48],pp21[47],pp22[46]},gpcOutL1_66);
wire [2:0] gpcOutL1_67;

// (* RLOC = "X1Y67" *)
gpc006 gpcL1_67 ({pp17[57],pp18[56],pp19[55],pp20[54],pp21[53],pp22[52]},gpcOutL1_67);
wire [2:0] gpcOutL1_68;

// (* RLOC = "X1Y68" *)
gpc006 gpcL1_68 ({pp17[63],pp18[62],pp19[61],pp20[60],pp21[59],pp22[58]},gpcOutL1_68);
wire [2:0] gpcOutL1_69;

// (* RLOC = "X1Y69" *)
gpc006 gpcL1_69 ({pp0[45],pp1[44],pp2[43],pp3[42],pp4[41],pp5[40]},gpcOutL1_69);
wire [2:0] gpcOutL1_70;

// (* RLOC = "X1Y70" *)
gpc006 gpcL1_70 ({pp6[45],pp7[44],pp8[43],pp9[42],pp10[41],pp11[40]},gpcOutL1_70);
wire [2:0] gpcOutL1_71;

// (* RLOC = "X1Y71" *)
gpc006 gpcL1_71 ({pp12[45],pp13[44],pp14[43],pp15[42],pp16[41],pp17[40]},gpcOutL1_71);
wire [2:0] gpcOutL1_72;

// (* RLOC = "X1Y72" *)
gpc006 gpcL1_72 ({pp18[45],pp19[44],pp20[43],pp21[42],pp22[41],pp23[40]},gpcOutL1_72);
wire [2:0] gpcOutL1_73;

// (* RLOC = "X1Y73" *)
gpc006 gpcL1_73 ({pp18[51],pp19[50],pp20[49],pp21[48],pp22[47],pp23[46]},gpcOutL1_73);
wire [2:0] gpcOutL1_74;

// (* RLOC = "X1Y74" *)
gpc006 gpcL1_74 ({pp18[57],pp19[56],pp20[55],pp21[54],pp22[53],pp23[52]},gpcOutL1_74);
wire [2:0] gpcOutL1_75;

// (* RLOC = "X1Y75" *)
gpc006 gpcL1_75 ({pp18[63],pp19[62],pp20[61],pp21[60],pp22[59],pp23[58]},gpcOutL1_75);
wire [2:0] gpcOutL1_76;

// (* RLOC = "X1Y76" *)
gpc006 gpcL1_76 ({pp0[44],pp1[43],pp2[42],pp3[41],pp4[40],pp5[39]},gpcOutL1_76);
wire [2:0] gpcOutL1_77;

// (* RLOC = "X1Y77" *)
gpc006 gpcL1_77 ({pp6[44],pp7[43],pp8[42],pp9[41],pp10[40],pp11[39]},gpcOutL1_77);
wire [2:0] gpcOutL1_78;

// (* RLOC = "X1Y78" *)
gpc006 gpcL1_78 ({pp12[44],pp13[43],pp14[42],pp15[41],pp16[40],pp17[39]},gpcOutL1_78);
wire [2:0] gpcOutL1_79;

// (* RLOC = "X1Y79" *)
gpc006 gpcL1_79 ({pp18[44],pp19[43],pp20[42],pp21[41],pp22[40],pp23[39]},gpcOutL1_79);
wire [2:0] gpcOutL1_80;

// (* RLOC = "X1Y80" *)
gpc006 gpcL1_80 ({pp19[45],pp20[44],pp21[43],pp22[42],pp23[41],pp24[40]},gpcOutL1_80);
wire [2:0] gpcOutL1_81;

// (* RLOC = "X1Y81" *)
gpc006 gpcL1_81 ({pp19[51],pp20[50],pp21[49],pp22[48],pp23[47],pp24[46]},gpcOutL1_81);
wire [2:0] gpcOutL1_82;

// (* RLOC = "X1Y82" *)
gpc006 gpcL1_82 ({pp19[57],pp20[56],pp21[55],pp22[54],pp23[53],pp24[52]},gpcOutL1_82);
wire [2:0] gpcOutL1_83;

// (* RLOC = "X1Y83" *)
gpc006 gpcL1_83 ({pp19[63],pp20[62],pp21[61],pp22[60],pp23[59],pp24[58]},gpcOutL1_83);
wire [2:0] gpcOutL1_84;

// (* RLOC = "X1Y84" *)
gpc006 gpcL1_84 ({pp0[43],pp1[42],pp2[41],pp3[40],pp4[39],pp5[38]},gpcOutL1_84);
wire [2:0] gpcOutL1_85;

// (* RLOC = "X1Y85" *)
gpc006 gpcL1_85 ({pp6[43],pp7[42],pp8[41],pp9[40],pp10[39],pp11[38]},gpcOutL1_85);
wire [2:0] gpcOutL1_86;

// (* RLOC = "X1Y86" *)
gpc006 gpcL1_86 ({pp12[43],pp13[42],pp14[41],pp15[40],pp16[39],pp17[38]},gpcOutL1_86);
wire [2:0] gpcOutL1_87;

// (* RLOC = "X1Y87" *)
gpc006 gpcL1_87 ({pp18[43],pp19[42],pp20[41],pp21[40],pp22[39],pp23[38]},gpcOutL1_87);
wire [2:0] gpcOutL1_88;

// (* RLOC = "X1Y88" *)
gpc006 gpcL1_88 ({pp20[45],pp21[44],pp22[43],pp23[42],pp24[41],pp25[40]},gpcOutL1_88);
wire [2:0] gpcOutL1_89;

// (* RLOC = "X1Y89" *)
gpc006 gpcL1_89 ({pp20[51],pp21[50],pp22[49],pp23[48],pp24[47],pp25[46]},gpcOutL1_89);
wire [2:0] gpcOutL1_90;

// (* RLOC = "X1Y90" *)
gpc006 gpcL1_90 ({pp20[57],pp21[56],pp22[55],pp23[54],pp24[53],pp25[52]},gpcOutL1_90);
wire [2:0] gpcOutL1_91;

// (* RLOC = "X1Y91" *)
gpc006 gpcL1_91 ({pp20[63],pp21[62],pp22[61],pp23[60],pp24[59],pp25[58]},gpcOutL1_91);
wire [2:0] gpcOutL1_92;

// (* RLOC = "X1Y92" *)
gpc006 gpcL1_92 ({pp0[42],pp1[41],pp2[40],pp3[39],pp4[38],pp5[37]},gpcOutL1_92);
wire [2:0] gpcOutL1_93;

// (* RLOC = "X1Y93" *)
gpc006 gpcL1_93 ({pp6[42],pp7[41],pp8[40],pp9[39],pp10[38],pp11[37]},gpcOutL1_93);
wire [2:0] gpcOutL1_94;

// (* RLOC = "X1Y94" *)
gpc006 gpcL1_94 ({pp12[42],pp13[41],pp14[40],pp15[39],pp16[38],pp17[37]},gpcOutL1_94);
wire [2:0] gpcOutL1_95;

// (* RLOC = "X1Y95" *)
gpc006 gpcL1_95 ({pp18[42],pp19[41],pp20[40],pp21[39],pp22[38],pp23[37]},gpcOutL1_95);
wire [2:0] gpcOutL1_96;

// (* RLOC = "X1Y96" *)
gpc006 gpcL1_96 ({pp21[45],pp22[44],pp23[43],pp24[42],pp25[41],pp26[40]},gpcOutL1_96);
wire [2:0] gpcOutL1_97;

// (* RLOC = "X1Y97" *)
gpc006 gpcL1_97 ({pp21[51],pp22[50],pp23[49],pp24[48],pp25[47],pp26[46]},gpcOutL1_97);
wire [2:0] gpcOutL1_98;

// (* RLOC = "X1Y98" *)
gpc006 gpcL1_98 ({pp21[57],pp22[56],pp23[55],pp24[54],pp25[53],pp26[52]},gpcOutL1_98);
wire [2:0] gpcOutL1_99;

// (* RLOC = "X1Y99" *)
gpc006 gpcL1_99 ({pp21[63],pp22[62],pp23[61],pp24[60],pp25[59],pp26[58]},gpcOutL1_99);
wire [2:0] gpcOutL1_100;

// (* RLOC = "X1Y100" *)
gpc006 gpcL1_100 ({pp0[41],pp1[40],pp2[39],pp3[38],pp4[37],pp5[36]},gpcOutL1_100);
wire [2:0] gpcOutL1_101;

// (* RLOC = "X1Y101" *)
gpc006 gpcL1_101 ({pp6[41],pp7[40],pp8[39],pp9[38],pp10[37],pp11[36]},gpcOutL1_101);
wire [2:0] gpcOutL1_102;

// (* RLOC = "X1Y102" *)
gpc006 gpcL1_102 ({pp12[41],pp13[40],pp14[39],pp15[38],pp16[37],pp17[36]},gpcOutL1_102);
wire [2:0] gpcOutL1_103;

// (* RLOC = "X1Y103" *)
gpc006 gpcL1_103 ({pp18[41],pp19[40],pp20[39],pp21[38],pp22[37],pp23[36]},gpcOutL1_103);
wire [2:0] gpcOutL1_104;

// (* RLOC = "X1Y104" *)
gpc006 gpcL1_104 ({pp22[45],pp23[44],pp24[43],pp25[42],pp26[41],pp27[40]},gpcOutL1_104);
wire [2:0] gpcOutL1_105;

// (* RLOC = "X1Y105" *)
gpc006 gpcL1_105 ({pp22[51],pp23[50],pp24[49],pp25[48],pp26[47],pp27[46]},gpcOutL1_105);
wire [2:0] gpcOutL1_106;

// (* RLOC = "X1Y106" *)
gpc006 gpcL1_106 ({pp22[57],pp23[56],pp24[55],pp25[54],pp26[53],pp27[52]},gpcOutL1_106);
wire [2:0] gpcOutL1_107;

// (* RLOC = "X1Y107" *)
gpc006 gpcL1_107 ({pp22[63],pp23[62],pp24[61],pp25[60],pp26[59],pp27[58]},gpcOutL1_107);
wire [2:0] gpcOutL1_108;

// (* RLOC = "X1Y108" *)
gpc006 gpcL1_108 ({pp0[40],pp1[39],pp2[38],pp3[37],pp4[36],pp5[35]},gpcOutL1_108);
wire [2:0] gpcOutL1_109;

// (* RLOC = "X1Y109" *)
gpc006 gpcL1_109 ({pp6[40],pp7[39],pp8[38],pp9[37],pp10[36],pp11[35]},gpcOutL1_109);
wire [2:0] gpcOutL1_110;

// (* RLOC = "X1Y110" *)
gpc006 gpcL1_110 ({pp12[40],pp13[39],pp14[38],pp15[37],pp16[36],pp17[35]},gpcOutL1_110);
wire [2:0] gpcOutL1_111;

// (* RLOC = "X1Y111" *)
gpc006 gpcL1_111 ({pp18[40],pp19[39],pp20[38],pp21[37],pp22[36],pp23[35]},gpcOutL1_111);
wire [2:0] gpcOutL1_112;

// (* RLOC = "X1Y112" *)
gpc006 gpcL1_112 ({pp23[45],pp24[44],pp25[43],pp26[42],pp27[41],pp28[40]},gpcOutL1_112);
wire [2:0] gpcOutL1_113;

// (* RLOC = "X1Y113" *)
gpc006 gpcL1_113 ({pp23[51],pp24[50],pp25[49],pp26[48],pp27[47],pp28[46]},gpcOutL1_113);
wire [2:0] gpcOutL1_114;

// (* RLOC = "X1Y114" *)
gpc006 gpcL1_114 ({pp23[57],pp24[56],pp25[55],pp26[54],pp27[53],pp28[52]},gpcOutL1_114);
wire [2:0] gpcOutL1_115;

// (* RLOC = "X1Y115" *)
gpc006 gpcL1_115 ({pp23[63],pp24[62],pp25[61],pp26[60],pp27[59],pp28[58]},gpcOutL1_115);
wire [2:0] gpcOutL1_116;

// (* RLOC = "X1Y116" *)
gpc006 gpcL1_116 ({pp0[39],pp1[38],pp2[37],pp3[36],pp4[35],pp5[34]},gpcOutL1_116);
wire [2:0] gpcOutL1_117;

// (* RLOC = "X1Y117" *)
gpc006 gpcL1_117 ({pp6[39],pp7[38],pp8[37],pp9[36],pp10[35],pp11[34]},gpcOutL1_117);
wire [2:0] gpcOutL1_118;

// (* RLOC = "X1Y118" *)
gpc006 gpcL1_118 ({pp12[39],pp13[38],pp14[37],pp15[36],pp16[35],pp17[34]},gpcOutL1_118);
wire [2:0] gpcOutL1_119;

// (* RLOC = "X1Y119" *)
gpc006 gpcL1_119 ({pp18[39],pp19[38],pp20[37],pp21[36],pp22[35],pp23[34]},gpcOutL1_119);
wire [2:0] gpcOutL1_120;

// (* RLOC = "X1Y120" *)
gpc006 gpcL1_120 ({pp24[39],pp25[38],pp26[37],pp27[36],pp28[35],pp29[34]},gpcOutL1_120);
wire [2:0] gpcOutL1_121;

// (* RLOC = "X1Y121" *)
gpc006 gpcL1_121 ({pp24[45],pp25[44],pp26[43],pp27[42],pp28[41],pp29[40]},gpcOutL1_121);
wire [2:0] gpcOutL1_122;

// (* RLOC = "X1Y122" *)
gpc006 gpcL1_122 ({pp24[51],pp25[50],pp26[49],pp27[48],pp28[47],pp29[46]},gpcOutL1_122);
wire [2:0] gpcOutL1_123;

// (* RLOC = "X1Y123" *)
gpc006 gpcL1_123 ({pp24[57],pp25[56],pp26[55],pp27[54],pp28[53],pp29[52]},gpcOutL1_123);
wire [2:0] gpcOutL1_124;

// (* RLOC = "X1Y124" *)
gpc006 gpcL1_124 ({pp24[63],pp25[62],pp26[61],pp27[60],pp28[59],pp29[58]},gpcOutL1_124);
wire [2:0] gpcOutL1_125;

// (* RLOC = "X1Y125" *)
gpc006 gpcL1_125 ({pp0[38],pp1[37],pp2[36],pp3[35],pp4[34],pp5[33]},gpcOutL1_125);
wire [2:0] gpcOutL1_126;

// (* RLOC = "X1Y126" *)
gpc006 gpcL1_126 ({pp6[38],pp7[37],pp8[36],pp9[35],pp10[34],pp11[33]},gpcOutL1_126);
wire [2:0] gpcOutL1_127;

// (* RLOC = "X1Y127" *)
gpc006 gpcL1_127 ({pp12[38],pp13[37],pp14[36],pp15[35],pp16[34],pp17[33]},gpcOutL1_127);
wire [2:0] gpcOutL1_128;

// (* RLOC = "X1Y128" *)
gpc006 gpcL1_128 ({pp18[38],pp19[37],pp20[36],pp21[35],pp22[34],pp23[33]},gpcOutL1_128);
wire [2:0] gpcOutL1_129;

// (* RLOC = "X1Y129" *)
gpc006 gpcL1_129 ({pp24[38],pp25[37],pp26[36],pp27[35],pp28[34],pp29[33]},gpcOutL1_129);
wire [2:0] gpcOutL1_130;

// (* RLOC = "X1Y130" *)
gpc006 gpcL1_130 ({pp25[39],pp26[38],pp27[37],pp28[36],pp29[35],pp30[34]},gpcOutL1_130);
wire [2:0] gpcOutL1_131;

// (* RLOC = "X1Y131" *)
gpc006 gpcL1_131 ({pp25[45],pp26[44],pp27[43],pp28[42],pp29[41],pp30[40]},gpcOutL1_131);
wire [2:0] gpcOutL1_132;

// (* RLOC = "X1Y132" *)
gpc006 gpcL1_132 ({pp25[51],pp26[50],pp27[49],pp28[48],pp29[47],pp30[46]},gpcOutL1_132);
wire [2:0] gpcOutL1_133;

// (* RLOC = "X1Y133" *)
gpc006 gpcL1_133 ({pp25[57],pp26[56],pp27[55],pp28[54],pp29[53],pp30[52]},gpcOutL1_133);
wire [2:0] gpcOutL1_134;

// (* RLOC = "X1Y134" *)
gpc006 gpcL1_134 ({pp25[63],pp26[62],pp27[61],pp28[60],pp29[59],pp30[58]},gpcOutL1_134);
wire [2:0] gpcOutL1_135;

// (* RLOC = "X1Y135" *)
gpc006 gpcL1_135 ({pp0[37],pp1[36],pp2[35],pp3[34],pp4[33],pp5[32]},gpcOutL1_135);
wire [2:0] gpcOutL1_136;

// (* RLOC = "X1Y136" *)
gpc006 gpcL1_136 ({pp6[37],pp7[36],pp8[35],pp9[34],pp10[33],pp11[32]},gpcOutL1_136);
wire [2:0] gpcOutL1_137;

// (* RLOC = "X1Y137" *)
gpc006 gpcL1_137 ({pp12[37],pp13[36],pp14[35],pp15[34],pp16[33],pp17[32]},gpcOutL1_137);
wire [2:0] gpcOutL1_138;

// (* RLOC = "X1Y138" *)
gpc006 gpcL1_138 ({pp18[37],pp19[36],pp20[35],pp21[34],pp22[33],pp23[32]},gpcOutL1_138);
wire [2:0] gpcOutL1_139;

// (* RLOC = "X1Y139" *)
gpc006 gpcL1_139 ({pp24[37],pp25[36],pp26[35],pp27[34],pp28[33],pp29[32]},gpcOutL1_139);
wire [2:0] gpcOutL1_140;

// (* RLOC = "X1Y140" *)
gpc006 gpcL1_140 ({pp26[39],pp27[38],pp28[37],pp29[36],pp30[35],pp31[34]},gpcOutL1_140);
wire [2:0] gpcOutL1_141;

// (* RLOC = "X1Y141" *)
gpc006 gpcL1_141 ({pp26[45],pp27[44],pp28[43],pp29[42],pp30[41],pp31[40]},gpcOutL1_141);
wire [2:0] gpcOutL1_142;

// (* RLOC = "X1Y142" *)
gpc006 gpcL1_142 ({pp26[51],pp27[50],pp28[49],pp29[48],pp30[47],pp31[46]},gpcOutL1_142);
wire [2:0] gpcOutL1_143;

// (* RLOC = "X1Y143" *)
gpc006 gpcL1_143 ({pp26[57],pp27[56],pp28[55],pp29[54],pp30[53],pp31[52]},gpcOutL1_143);
wire [2:0] gpcOutL1_144;

// (* RLOC = "X1Y144" *)
gpc006 gpcL1_144 ({pp26[63],pp27[62],pp28[61],pp29[60],pp30[59],pp31[58]},gpcOutL1_144);
wire [2:0] gpcOutL1_145;

// (* RLOC = "X1Y145" *)
gpc006 gpcL1_145 ({pp0[36],pp1[35],pp2[34],pp3[33],pp4[32],pp5[31]},gpcOutL1_145);
wire [2:0] gpcOutL1_146;

// (* RLOC = "X1Y146" *)
gpc006 gpcL1_146 ({pp6[36],pp7[35],pp8[34],pp9[33],pp10[32],pp11[31]},gpcOutL1_146);
wire [2:0] gpcOutL1_147;

// (* RLOC = "X1Y147" *)
gpc006 gpcL1_147 ({pp12[36],pp13[35],pp14[34],pp15[33],pp16[32],pp17[31]},gpcOutL1_147);
wire [2:0] gpcOutL1_148;

// (* RLOC = "X1Y148" *)
gpc006 gpcL1_148 ({pp18[36],pp19[35],pp20[34],pp21[33],pp22[32],pp23[31]},gpcOutL1_148);
wire [2:0] gpcOutL1_149;

// (* RLOC = "X1Y149" *)
gpc006 gpcL1_149 ({pp24[36],pp25[35],pp26[34],pp27[33],pp28[32],pp29[31]},gpcOutL1_149);
wire [2:0] gpcOutL1_150;

// (* RLOC = "X1Y150" *)
gpc006 gpcL1_150 ({pp27[39],pp28[38],pp29[37],pp30[36],pp31[35],pp32[34]},gpcOutL1_150);
wire [2:0] gpcOutL1_151;

// (* RLOC = "X1Y151" *)
gpc006 gpcL1_151 ({pp27[45],pp28[44],pp29[43],pp30[42],pp31[41],pp32[40]},gpcOutL1_151);
wire [2:0] gpcOutL1_152;

// (* RLOC = "X1Y152" *)
gpc006 gpcL1_152 ({pp27[51],pp28[50],pp29[49],pp30[48],pp31[47],pp32[46]},gpcOutL1_152);
wire [2:0] gpcOutL1_153;

// (* RLOC = "X1Y153" *)
gpc006 gpcL1_153 ({pp27[57],pp28[56],pp29[55],pp30[54],pp31[53],pp32[52]},gpcOutL1_153);
wire [2:0] gpcOutL1_154;

// (* RLOC = "X1Y154" *)
gpc006 gpcL1_154 ({pp27[63],pp28[62],pp29[61],pp30[60],pp31[59],pp32[58]},gpcOutL1_154);
wire [2:0] gpcOutL1_155;

// (* RLOC = "X1Y155" *)
gpc006 gpcL1_155 ({pp0[35],pp1[34],pp2[33],pp3[32],pp4[31],pp5[30]},gpcOutL1_155);
wire [2:0] gpcOutL1_156;

// (* RLOC = "X1Y156" *)
gpc006 gpcL1_156 ({pp6[35],pp7[34],pp8[33],pp9[32],pp10[31],pp11[30]},gpcOutL1_156);
wire [2:0] gpcOutL1_157;

// (* RLOC = "X1Y157" *)
gpc006 gpcL1_157 ({pp12[35],pp13[34],pp14[33],pp15[32],pp16[31],pp17[30]},gpcOutL1_157);
wire [2:0] gpcOutL1_158;

// (* RLOC = "X1Y158" *)
gpc006 gpcL1_158 ({pp18[35],pp19[34],pp20[33],pp21[32],pp22[31],pp23[30]},gpcOutL1_158);
wire [2:0] gpcOutL1_159;

// (* RLOC = "X1Y159" *)
gpc006 gpcL1_159 ({pp24[35],pp25[34],pp26[33],pp27[32],pp28[31],pp29[30]},gpcOutL1_159);
wire [2:0] gpcOutL1_160;

// (* RLOC = "X1Y160" *)
gpc006 gpcL1_160 ({pp28[39],pp29[38],pp30[37],pp31[36],pp32[35],pp33[34]},gpcOutL1_160);
wire [2:0] gpcOutL1_161;

// (* RLOC = "X1Y161" *)
gpc006 gpcL1_161 ({pp28[45],pp29[44],pp30[43],pp31[42],pp32[41],pp33[40]},gpcOutL1_161);
wire [2:0] gpcOutL1_162;

// (* RLOC = "X1Y162" *)
gpc006 gpcL1_162 ({pp28[51],pp29[50],pp30[49],pp31[48],pp32[47],pp33[46]},gpcOutL1_162);
wire [2:0] gpcOutL1_163;

// (* RLOC = "X1Y163" *)
gpc006 gpcL1_163 ({pp28[57],pp29[56],pp30[55],pp31[54],pp32[53],pp33[52]},gpcOutL1_163);
wire [2:0] gpcOutL1_164;

// (* RLOC = "X1Y164" *)
gpc006 gpcL1_164 ({pp28[63],pp29[62],pp30[61],pp31[60],pp32[59],pp33[58]},gpcOutL1_164);
wire [2:0] gpcOutL1_165;

// (* RLOC = "X1Y165" *)
gpc006 gpcL1_165 ({pp0[34],pp1[33],pp2[32],pp3[31],pp4[30],pp5[29]},gpcOutL1_165);
wire [2:0] gpcOutL1_166;

// (* RLOC = "X1Y166" *)
gpc006 gpcL1_166 ({pp6[34],pp7[33],pp8[32],pp9[31],pp10[30],pp11[29]},gpcOutL1_166);
wire [2:0] gpcOutL1_167;

// (* RLOC = "X1Y167" *)
gpc006 gpcL1_167 ({pp12[34],pp13[33],pp14[32],pp15[31],pp16[30],pp17[29]},gpcOutL1_167);
wire [2:0] gpcOutL1_168;

// (* RLOC = "X1Y168" *)
gpc006 gpcL1_168 ({pp18[34],pp19[33],pp20[32],pp21[31],pp22[30],pp23[29]},gpcOutL1_168);
wire [2:0] gpcOutL1_169;

// (* RLOC = "X1Y169" *)
gpc006 gpcL1_169 ({pp24[34],pp25[33],pp26[32],pp27[31],pp28[30],pp29[29]},gpcOutL1_169);
wire [2:0] gpcOutL1_170;

// (* RLOC = "X1Y170" *)
gpc006 gpcL1_170 ({pp29[39],pp30[38],pp31[37],pp32[36],pp33[35],pp34[34]},gpcOutL1_170);
wire [2:0] gpcOutL1_171;

// (* RLOC = "X1Y171" *)
gpc006 gpcL1_171 ({pp29[45],pp30[44],pp31[43],pp32[42],pp33[41],pp34[40]},gpcOutL1_171);
wire [2:0] gpcOutL1_172;

// (* RLOC = "X1Y172" *)
gpc006 gpcL1_172 ({pp29[51],pp30[50],pp31[49],pp32[48],pp33[47],pp34[46]},gpcOutL1_172);
wire [2:0] gpcOutL1_173;

// (* RLOC = "X1Y173" *)
gpc006 gpcL1_173 ({pp29[57],pp30[56],pp31[55],pp32[54],pp33[53],pp34[52]},gpcOutL1_173);
wire [2:0] gpcOutL1_174;

// (* RLOC = "X1Y174" *)
gpc006 gpcL1_174 ({pp29[63],pp30[62],pp31[61],pp32[60],pp33[59],pp34[58]},gpcOutL1_174);
wire [2:0] gpcOutL1_175;

// (* RLOC = "X1Y175" *)
gpc006 gpcL1_175 ({pp0[33],pp1[32],pp2[31],pp3[30],pp4[29],pp5[28]},gpcOutL1_175);
wire [2:0] gpcOutL1_176;

// (* RLOC = "X1Y176" *)
gpc006 gpcL1_176 ({pp6[33],pp7[32],pp8[31],pp9[30],pp10[29],pp11[28]},gpcOutL1_176);
wire [2:0] gpcOutL1_177;

// (* RLOC = "X1Y177" *)
gpc006 gpcL1_177 ({pp12[33],pp13[32],pp14[31],pp15[30],pp16[29],pp17[28]},gpcOutL1_177);
wire [2:0] gpcOutL1_178;

// (* RLOC = "X1Y178" *)
gpc006 gpcL1_178 ({pp18[33],pp19[32],pp20[31],pp21[30],pp22[29],pp23[28]},gpcOutL1_178);
wire [2:0] gpcOutL1_179;

// (* RLOC = "X1Y179" *)
gpc006 gpcL1_179 ({pp24[33],pp25[32],pp26[31],pp27[30],pp28[29],pp29[28]},gpcOutL1_179);
wire [2:0] gpcOutL1_180;

// (* RLOC = "X1Y180" *)
gpc006 gpcL1_180 ({pp30[33],pp31[32],pp32[31],pp33[30],pp34[29],pp35[28]},gpcOutL1_180);
wire [2:0] gpcOutL1_181;

// (* RLOC = "X1Y181" *)
gpc006 gpcL1_181 ({pp30[39],pp31[38],pp32[37],pp33[36],pp34[35],pp35[34]},gpcOutL1_181);
wire [2:0] gpcOutL1_182;

// (* RLOC = "X1Y182" *)
gpc006 gpcL1_182 ({pp30[45],pp31[44],pp32[43],pp33[42],pp34[41],pp35[40]},gpcOutL1_182);
wire [2:0] gpcOutL1_183;

// (* RLOC = "X1Y183" *)
gpc006 gpcL1_183 ({pp30[51],pp31[50],pp32[49],pp33[48],pp34[47],pp35[46]},gpcOutL1_183);
wire [2:0] gpcOutL1_184;

// (* RLOC = "X1Y184" *)
gpc006 gpcL1_184 ({pp30[57],pp31[56],pp32[55],pp33[54],pp34[53],pp35[52]},gpcOutL1_184);
wire [2:0] gpcOutL1_185;

// (* RLOC = "X1Y185" *)
gpc006 gpcL1_185 ({pp30[63],pp31[62],pp32[61],pp33[60],pp34[59],pp35[58]},gpcOutL1_185);
wire [2:0] gpcOutL1_186;

// (* RLOC = "X1Y186" *)
gpc006 gpcL1_186 ({pp0[32],pp1[31],pp2[30],pp3[29],pp4[28],pp5[27]},gpcOutL1_186);
wire [2:0] gpcOutL1_187;

// (* RLOC = "X1Y187" *)
gpc006 gpcL1_187 ({pp6[32],pp7[31],pp8[30],pp9[29],pp10[28],pp11[27]},gpcOutL1_187);
wire [2:0] gpcOutL1_188;

// (* RLOC = "X1Y188" *)
gpc006 gpcL1_188 ({pp12[32],pp13[31],pp14[30],pp15[29],pp16[28],pp17[27]},gpcOutL1_188);
wire [2:0] gpcOutL1_189;

// (* RLOC = "X1Y189" *)
gpc006 gpcL1_189 ({pp18[32],pp19[31],pp20[30],pp21[29],pp22[28],pp23[27]},gpcOutL1_189);
wire [2:0] gpcOutL1_190;

// (* RLOC = "X1Y190" *)
gpc006 gpcL1_190 ({pp24[32],pp25[31],pp26[30],pp27[29],pp28[28],pp29[27]},gpcOutL1_190);
wire [2:0] gpcOutL1_191;

// (* RLOC = "X1Y191" *)
gpc006 gpcL1_191 ({pp30[32],pp31[31],pp32[30],pp33[29],pp34[28],pp35[27]},gpcOutL1_191);
wire [2:0] gpcOutL1_192;

// (* RLOC = "X1Y192" *)
gpc006 gpcL1_192 ({pp31[33],pp32[32],pp33[31],pp34[30],pp35[29],pp36[28]},gpcOutL1_192);
wire [2:0] gpcOutL1_193;

// (* RLOC = "X1Y193" *)
gpc006 gpcL1_193 ({pp31[39],pp32[38],pp33[37],pp34[36],pp35[35],pp36[34]},gpcOutL1_193);
wire [2:0] gpcOutL1_194;

// (* RLOC = "X1Y194" *)
gpc006 gpcL1_194 ({pp31[45],pp32[44],pp33[43],pp34[42],pp35[41],pp36[40]},gpcOutL1_194);
wire [2:0] gpcOutL1_195;

// (* RLOC = "X1Y195" *)
gpc006 gpcL1_195 ({pp31[51],pp32[50],pp33[49],pp34[48],pp35[47],pp36[46]},gpcOutL1_195);
wire [2:0] gpcOutL1_196;

// (* RLOC = "X1Y196" *)
gpc006 gpcL1_196 ({pp31[57],pp32[56],pp33[55],pp34[54],pp35[53],pp36[52]},gpcOutL1_196);
wire [2:0] gpcOutL1_197;

// (* RLOC = "X1Y197" *)
gpc006 gpcL1_197 ({pp31[63],pp32[62],pp33[61],pp34[60],pp35[59],pp36[58]},gpcOutL1_197);
wire [2:0] gpcOutL1_198;

// (* RLOC = "X1Y198" *)
gpc006 gpcL1_198 ({pp0[31],pp1[30],pp2[29],pp3[28],pp4[27],pp5[26]},gpcOutL1_198);
wire [2:0] gpcOutL1_199;

// (* RLOC = "X1Y199" *)
gpc006 gpcL1_199 ({pp6[31],pp7[30],pp8[29],pp9[28],pp10[27],pp11[26]},gpcOutL1_199);
wire [2:0] gpcOutL1_200;

// (* RLOC = "X1Y200" *)
gpc006 gpcL1_200 ({pp12[31],pp13[30],pp14[29],pp15[28],pp16[27],pp17[26]},gpcOutL1_200);
wire [2:0] gpcOutL1_201;

// (* RLOC = "X1Y201" *)
gpc006 gpcL1_201 ({pp18[31],pp19[30],pp20[29],pp21[28],pp22[27],pp23[26]},gpcOutL1_201);
wire [2:0] gpcOutL1_202;

// (* RLOC = "X1Y202" *)
gpc006 gpcL1_202 ({pp24[31],pp25[30],pp26[29],pp27[28],pp28[27],pp29[26]},gpcOutL1_202);
wire [2:0] gpcOutL1_203;

// (* RLOC = "X1Y203" *)
gpc006 gpcL1_203 ({pp30[31],pp31[30],pp32[29],pp33[28],pp34[27],pp35[26]},gpcOutL1_203);
wire [2:0] gpcOutL1_204;

// (* RLOC = "X1Y204" *)
gpc006 gpcL1_204 ({pp32[33],pp33[32],pp34[31],pp35[30],pp36[29],pp37[28]},gpcOutL1_204);
wire [2:0] gpcOutL1_205;

// (* RLOC = "X1Y205" *)
gpc006 gpcL1_205 ({pp32[39],pp33[38],pp34[37],pp35[36],pp36[35],pp37[34]},gpcOutL1_205);
wire [2:0] gpcOutL1_206;

// (* RLOC = "X1Y206" *)
gpc006 gpcL1_206 ({pp32[45],pp33[44],pp34[43],pp35[42],pp36[41],pp37[40]},gpcOutL1_206);
wire [2:0] gpcOutL1_207;

// (* RLOC = "X1Y207" *)
gpc006 gpcL1_207 ({pp32[51],pp33[50],pp34[49],pp35[48],pp36[47],pp37[46]},gpcOutL1_207);
wire [2:0] gpcOutL1_208;

// (* RLOC = "X1Y208" *)
gpc006 gpcL1_208 ({pp32[57],pp33[56],pp34[55],pp35[54],pp36[53],pp37[52]},gpcOutL1_208);
wire [2:0] gpcOutL1_209;

// (* RLOC = "X1Y209" *)
gpc006 gpcL1_209 ({pp32[63],pp33[62],pp34[61],pp35[60],pp36[59],pp37[58]},gpcOutL1_209);
wire [2:0] gpcOutL1_210;

// (* RLOC = "X1Y210" *)
gpc006 gpcL1_210 ({pp0[30],pp1[29],pp2[28],pp3[27],pp4[26],pp5[25]},gpcOutL1_210);
wire [2:0] gpcOutL1_211;

// (* RLOC = "X1Y211" *)
gpc006 gpcL1_211 ({pp6[30],pp7[29],pp8[28],pp9[27],pp10[26],pp11[25]},gpcOutL1_211);
wire [2:0] gpcOutL1_212;

// (* RLOC = "X1Y212" *)
gpc006 gpcL1_212 ({pp12[30],pp13[29],pp14[28],pp15[27],pp16[26],pp17[25]},gpcOutL1_212);
wire [2:0] gpcOutL1_213;

// (* RLOC = "X1Y213" *)
gpc006 gpcL1_213 ({pp18[30],pp19[29],pp20[28],pp21[27],pp22[26],pp23[25]},gpcOutL1_213);
wire [2:0] gpcOutL1_214;

// (* RLOC = "X1Y214" *)
gpc006 gpcL1_214 ({pp24[30],pp25[29],pp26[28],pp27[27],pp28[26],pp29[25]},gpcOutL1_214);
wire [2:0] gpcOutL1_215;

// (* RLOC = "X1Y215" *)
gpc006 gpcL1_215 ({pp30[30],pp31[29],pp32[28],pp33[27],pp34[26],pp35[25]},gpcOutL1_215);
wire [2:0] gpcOutL1_216;

// (* RLOC = "X1Y216" *)
gpc006 gpcL1_216 ({pp33[33],pp34[32],pp35[31],pp36[30],pp37[29],pp38[28]},gpcOutL1_216);
wire [2:0] gpcOutL1_217;

// (* RLOC = "X1Y217" *)
gpc006 gpcL1_217 ({pp33[39],pp34[38],pp35[37],pp36[36],pp37[35],pp38[34]},gpcOutL1_217);
wire [2:0] gpcOutL1_218;

// (* RLOC = "X1Y218" *)
gpc006 gpcL1_218 ({pp33[45],pp34[44],pp35[43],pp36[42],pp37[41],pp38[40]},gpcOutL1_218);
wire [2:0] gpcOutL1_219;

// (* RLOC = "X1Y219" *)
gpc006 gpcL1_219 ({pp33[51],pp34[50],pp35[49],pp36[48],pp37[47],pp38[46]},gpcOutL1_219);
wire [2:0] gpcOutL1_220;

// (* RLOC = "X1Y220" *)
gpc006 gpcL1_220 ({pp33[57],pp34[56],pp35[55],pp36[54],pp37[53],pp38[52]},gpcOutL1_220);
wire [2:0] gpcOutL1_221;

// (* RLOC = "X1Y221" *)
gpc006 gpcL1_221 ({pp33[63],pp34[62],pp35[61],pp36[60],pp37[59],pp38[58]},gpcOutL1_221);
wire [2:0] gpcOutL1_222;

// (* RLOC = "X1Y222" *)
gpc006 gpcL1_222 ({pp0[29],pp1[28],pp2[27],pp3[26],pp4[25],pp5[24]},gpcOutL1_222);
wire [2:0] gpcOutL1_223;

// (* RLOC = "X1Y223" *)
gpc006 gpcL1_223 ({pp6[29],pp7[28],pp8[27],pp9[26],pp10[25],pp11[24]},gpcOutL1_223);
wire [2:0] gpcOutL1_224;

// (* RLOC = "X1Y224" *)
gpc006 gpcL1_224 ({pp12[29],pp13[28],pp14[27],pp15[26],pp16[25],pp17[24]},gpcOutL1_224);
wire [2:0] gpcOutL1_225;

// (* RLOC = "X1Y225" *)
gpc006 gpcL1_225 ({pp18[29],pp19[28],pp20[27],pp21[26],pp22[25],pp23[24]},gpcOutL1_225);
wire [2:0] gpcOutL1_226;

// (* RLOC = "X1Y226" *)
gpc006 gpcL1_226 ({pp24[29],pp25[28],pp26[27],pp27[26],pp28[25],pp29[24]},gpcOutL1_226);
wire [2:0] gpcOutL1_227;

// (* RLOC = "X1Y227" *)
gpc006 gpcL1_227 ({pp30[29],pp31[28],pp32[27],pp33[26],pp34[25],pp35[24]},gpcOutL1_227);
wire [2:0] gpcOutL1_228;

// (* RLOC = "X1Y228" *)
gpc006 gpcL1_228 ({pp34[33],pp35[32],pp36[31],pp37[30],pp38[29],pp39[28]},gpcOutL1_228);
wire [2:0] gpcOutL1_229;

// (* RLOC = "X1Y229" *)
gpc006 gpcL1_229 ({pp34[39],pp35[38],pp36[37],pp37[36],pp38[35],pp39[34]},gpcOutL1_229);
wire [2:0] gpcOutL1_230;

// (* RLOC = "X1Y230" *)
gpc006 gpcL1_230 ({pp34[45],pp35[44],pp36[43],pp37[42],pp38[41],pp39[40]},gpcOutL1_230);
wire [2:0] gpcOutL1_231;

// (* RLOC = "X1Y231" *)
gpc006 gpcL1_231 ({pp34[51],pp35[50],pp36[49],pp37[48],pp38[47],pp39[46]},gpcOutL1_231);
wire [2:0] gpcOutL1_232;

// (* RLOC = "X1Y232" *)
gpc006 gpcL1_232 ({pp34[57],pp35[56],pp36[55],pp37[54],pp38[53],pp39[52]},gpcOutL1_232);
wire [2:0] gpcOutL1_233;

// (* RLOC = "X1Y233" *)
gpc006 gpcL1_233 ({pp34[63],pp35[62],pp36[61],pp37[60],pp38[59],pp39[58]},gpcOutL1_233);
wire [2:0] gpcOutL1_234;

// (* RLOC = "X1Y234" *)
gpc006 gpcL1_234 ({pp0[28],pp1[27],pp2[26],pp3[25],pp4[24],pp5[23]},gpcOutL1_234);
wire [2:0] gpcOutL1_235;

// (* RLOC = "X1Y235" *)
gpc006 gpcL1_235 ({pp6[28],pp7[27],pp8[26],pp9[25],pp10[24],pp11[23]},gpcOutL1_235);
wire [2:0] gpcOutL1_236;

// (* RLOC = "X1Y236" *)
gpc006 gpcL1_236 ({pp12[28],pp13[27],pp14[26],pp15[25],pp16[24],pp17[23]},gpcOutL1_236);
wire [2:0] gpcOutL1_237;

// (* RLOC = "X1Y237" *)
gpc006 gpcL1_237 ({pp18[28],pp19[27],pp20[26],pp21[25],pp22[24],pp23[23]},gpcOutL1_237);
wire [2:0] gpcOutL1_238;

// (* RLOC = "X1Y238" *)
gpc006 gpcL1_238 ({pp24[28],pp25[27],pp26[26],pp27[25],pp28[24],pp29[23]},gpcOutL1_238);
wire [2:0] gpcOutL1_239;

// (* RLOC = "X1Y239" *)
gpc006 gpcL1_239 ({pp30[28],pp31[27],pp32[26],pp33[25],pp34[24],pp35[23]},gpcOutL1_239);
wire [2:0] gpcOutL1_240;

// (* RLOC = "X1Y240" *)
gpc006 gpcL1_240 ({pp35[33],pp36[32],pp37[31],pp38[30],pp39[29],pp40[28]},gpcOutL1_240);
wire [2:0] gpcOutL1_241;

// (* RLOC = "X1Y241" *)
gpc006 gpcL1_241 ({pp35[39],pp36[38],pp37[37],pp38[36],pp39[35],pp40[34]},gpcOutL1_241);
wire [2:0] gpcOutL1_242;

// (* RLOC = "X1Y242" *)
gpc006 gpcL1_242 ({pp35[45],pp36[44],pp37[43],pp38[42],pp39[41],pp40[40]},gpcOutL1_242);
wire [2:0] gpcOutL1_243;

// (* RLOC = "X1Y243" *)
gpc006 gpcL1_243 ({pp35[51],pp36[50],pp37[49],pp38[48],pp39[47],pp40[46]},gpcOutL1_243);
wire [2:0] gpcOutL1_244;

// (* RLOC = "X1Y244" *)
gpc006 gpcL1_244 ({pp35[57],pp36[56],pp37[55],pp38[54],pp39[53],pp40[52]},gpcOutL1_244);
wire [2:0] gpcOutL1_245;

// (* RLOC = "X1Y245" *)
gpc006 gpcL1_245 ({pp35[63],pp36[62],pp37[61],pp38[60],pp39[59],pp40[58]},gpcOutL1_245);
wire [2:0] gpcOutL1_246;

// (* RLOC = "X1Y246" *)
gpc006 gpcL1_246 ({pp0[27],pp1[26],pp2[25],pp3[24],pp4[23],pp5[22]},gpcOutL1_246);
wire [2:0] gpcOutL1_247;

// (* RLOC = "X1Y247" *)
gpc006 gpcL1_247 ({pp6[27],pp7[26],pp8[25],pp9[24],pp10[23],pp11[22]},gpcOutL1_247);
wire [2:0] gpcOutL1_248;

// (* RLOC = "X1Y248" *)
gpc006 gpcL1_248 ({pp12[27],pp13[26],pp14[25],pp15[24],pp16[23],pp17[22]},gpcOutL1_248);
wire [2:0] gpcOutL1_249;

// (* RLOC = "X1Y249" *)
gpc006 gpcL1_249 ({pp18[27],pp19[26],pp20[25],pp21[24],pp22[23],pp23[22]},gpcOutL1_249);
wire [2:0] gpcOutL1_250;

// (* RLOC = "X1Y250" *)
gpc006 gpcL1_250 ({pp24[27],pp25[26],pp26[25],pp27[24],pp28[23],pp29[22]},gpcOutL1_250);
wire [2:0] gpcOutL1_251;

// (* RLOC = "X1Y251" *)
gpc006 gpcL1_251 ({pp30[27],pp31[26],pp32[25],pp33[24],pp34[23],pp35[22]},gpcOutL1_251);
wire [2:0] gpcOutL1_252;

// (* RLOC = "X1Y252" *)
gpc006 gpcL1_252 ({pp36[27],pp37[26],pp38[25],pp39[24],pp40[23],pp41[22]},gpcOutL1_252);
wire [2:0] gpcOutL1_253;

// (* RLOC = "X1Y253" *)
gpc006 gpcL1_253 ({pp36[33],pp37[32],pp38[31],pp39[30],pp40[29],pp41[28]},gpcOutL1_253);
wire [2:0] gpcOutL1_254;

// (* RLOC = "X1Y254" *)
gpc006 gpcL1_254 ({pp36[39],pp37[38],pp38[37],pp39[36],pp40[35],pp41[34]},gpcOutL1_254);
wire [2:0] gpcOutL1_255;

// (* RLOC = "X1Y255" *)
gpc006 gpcL1_255 ({pp36[45],pp37[44],pp38[43],pp39[42],pp40[41],pp41[40]},gpcOutL1_255);
wire [2:0] gpcOutL1_256;

// (* RLOC = "X1Y256" *)
gpc006 gpcL1_256 ({pp36[51],pp37[50],pp38[49],pp39[48],pp40[47],pp41[46]},gpcOutL1_256);
wire [2:0] gpcOutL1_257;

// (* RLOC = "X1Y257" *)
gpc006 gpcL1_257 ({pp36[57],pp37[56],pp38[55],pp39[54],pp40[53],pp41[52]},gpcOutL1_257);
wire [2:0] gpcOutL1_258;

// (* RLOC = "X1Y258" *)
gpc006 gpcL1_258 ({pp36[63],pp37[62],pp38[61],pp39[60],pp40[59],pp41[58]},gpcOutL1_258);
wire [2:0] gpcOutL1_259;

// (* RLOC = "X1Y259" *)
gpc006 gpcL1_259 ({pp0[26],pp1[25],pp2[24],pp3[23],pp4[22],pp5[21]},gpcOutL1_259);
wire [2:0] gpcOutL1_260;

// (* RLOC = "X1Y260" *)
gpc006 gpcL1_260 ({pp6[26],pp7[25],pp8[24],pp9[23],pp10[22],pp11[21]},gpcOutL1_260);
wire [2:0] gpcOutL1_261;

// (* RLOC = "X1Y261" *)
gpc006 gpcL1_261 ({pp12[26],pp13[25],pp14[24],pp15[23],pp16[22],pp17[21]},gpcOutL1_261);
wire [2:0] gpcOutL1_262;

// (* RLOC = "X1Y262" *)
gpc006 gpcL1_262 ({pp18[26],pp19[25],pp20[24],pp21[23],pp22[22],pp23[21]},gpcOutL1_262);
wire [2:0] gpcOutL1_263;

// (* RLOC = "X1Y263" *)
gpc006 gpcL1_263 ({pp24[26],pp25[25],pp26[24],pp27[23],pp28[22],pp29[21]},gpcOutL1_263);
wire [2:0] gpcOutL1_264;

// (* RLOC = "X1Y264" *)
gpc006 gpcL1_264 ({pp30[26],pp31[25],pp32[24],pp33[23],pp34[22],pp35[21]},gpcOutL1_264);
wire [2:0] gpcOutL1_265;

// (* RLOC = "X1Y265" *)
gpc006 gpcL1_265 ({pp36[26],pp37[25],pp38[24],pp39[23],pp40[22],pp41[21]},gpcOutL1_265);
wire [2:0] gpcOutL1_266;

// (* RLOC = "X1Y266" *)
gpc006 gpcL1_266 ({pp37[27],pp38[26],pp39[25],pp40[24],pp41[23],pp42[22]},gpcOutL1_266);
wire [2:0] gpcOutL1_267;

// (* RLOC = "X1Y267" *)
gpc006 gpcL1_267 ({pp37[33],pp38[32],pp39[31],pp40[30],pp41[29],pp42[28]},gpcOutL1_267);
wire [2:0] gpcOutL1_268;

// (* RLOC = "X1Y268" *)
gpc006 gpcL1_268 ({pp37[39],pp38[38],pp39[37],pp40[36],pp41[35],pp42[34]},gpcOutL1_268);
wire [2:0] gpcOutL1_269;

// (* RLOC = "X1Y269" *)
gpc006 gpcL1_269 ({pp37[45],pp38[44],pp39[43],pp40[42],pp41[41],pp42[40]},gpcOutL1_269);
wire [2:0] gpcOutL1_270;

// (* RLOC = "X1Y270" *)
gpc006 gpcL1_270 ({pp37[51],pp38[50],pp39[49],pp40[48],pp41[47],pp42[46]},gpcOutL1_270);
wire [2:0] gpcOutL1_271;

// (* RLOC = "X1Y271" *)
gpc006 gpcL1_271 ({pp37[57],pp38[56],pp39[55],pp40[54],pp41[53],pp42[52]},gpcOutL1_271);
wire [2:0] gpcOutL1_272;

// (* RLOC = "X1Y272" *)
gpc006 gpcL1_272 ({pp37[63],pp38[62],pp39[61],pp40[60],pp41[59],pp42[58]},gpcOutL1_272);
wire [2:0] gpcOutL1_273;

// (* RLOC = "X1Y273" *)
gpc006 gpcL1_273 ({pp0[25],pp1[24],pp2[23],pp3[22],pp4[21],pp5[20]},gpcOutL1_273);
wire [2:0] gpcOutL1_274;

// (* RLOC = "X1Y274" *)
gpc006 gpcL1_274 ({pp6[25],pp7[24],pp8[23],pp9[22],pp10[21],pp11[20]},gpcOutL1_274);
wire [2:0] gpcOutL1_275;

// (* RLOC = "X1Y275" *)
gpc006 gpcL1_275 ({pp12[25],pp13[24],pp14[23],pp15[22],pp16[21],pp17[20]},gpcOutL1_275);
wire [2:0] gpcOutL1_276;

// (* RLOC = "X1Y276" *)
gpc006 gpcL1_276 ({pp18[25],pp19[24],pp20[23],pp21[22],pp22[21],pp23[20]},gpcOutL1_276);
wire [2:0] gpcOutL1_277;

// (* RLOC = "X1Y277" *)
gpc006 gpcL1_277 ({pp24[25],pp25[24],pp26[23],pp27[22],pp28[21],pp29[20]},gpcOutL1_277);
wire [2:0] gpcOutL1_278;

// (* RLOC = "X1Y278" *)
gpc006 gpcL1_278 ({pp30[25],pp31[24],pp32[23],pp33[22],pp34[21],pp35[20]},gpcOutL1_278);
wire [2:0] gpcOutL1_279;

// (* RLOC = "X1Y279" *)
gpc006 gpcL1_279 ({pp36[25],pp37[24],pp38[23],pp39[22],pp40[21],pp41[20]},gpcOutL1_279);
wire [2:0] gpcOutL1_280;

// (* RLOC = "X1Y280" *)
gpc006 gpcL1_280 ({pp38[27],pp39[26],pp40[25],pp41[24],pp42[23],pp43[22]},gpcOutL1_280);
wire [2:0] gpcOutL1_281;

// (* RLOC = "X1Y281" *)
gpc006 gpcL1_281 ({pp38[33],pp39[32],pp40[31],pp41[30],pp42[29],pp43[28]},gpcOutL1_281);
wire [2:0] gpcOutL1_282;

// (* RLOC = "X1Y282" *)
gpc006 gpcL1_282 ({pp38[39],pp39[38],pp40[37],pp41[36],pp42[35],pp43[34]},gpcOutL1_282);
wire [2:0] gpcOutL1_283;

// (* RLOC = "X1Y283" *)
gpc006 gpcL1_283 ({pp38[45],pp39[44],pp40[43],pp41[42],pp42[41],pp43[40]},gpcOutL1_283);
wire [2:0] gpcOutL1_284;

// (* RLOC = "X1Y284" *)
gpc006 gpcL1_284 ({pp38[51],pp39[50],pp40[49],pp41[48],pp42[47],pp43[46]},gpcOutL1_284);
wire [2:0] gpcOutL1_285;

// (* RLOC = "X1Y285" *)
gpc006 gpcL1_285 ({pp38[57],pp39[56],pp40[55],pp41[54],pp42[53],pp43[52]},gpcOutL1_285);
wire [2:0] gpcOutL1_286;

// (* RLOC = "X1Y286" *)
gpc006 gpcL1_286 ({pp38[63],pp39[62],pp40[61],pp41[60],pp42[59],pp43[58]},gpcOutL1_286);
wire [2:0] gpcOutL1_287;

// (* RLOC = "X1Y287" *)
gpc006 gpcL1_287 ({pp0[24],pp1[23],pp2[22],pp3[21],pp4[20],pp5[19]},gpcOutL1_287);
wire [2:0] gpcOutL1_288;

// (* RLOC = "X1Y288" *)
gpc006 gpcL1_288 ({pp6[24],pp7[23],pp8[22],pp9[21],pp10[20],pp11[19]},gpcOutL1_288);
wire [2:0] gpcOutL1_289;

// (* RLOC = "X1Y289" *)
gpc006 gpcL1_289 ({pp12[24],pp13[23],pp14[22],pp15[21],pp16[20],pp17[19]},gpcOutL1_289);
wire [2:0] gpcOutL1_290;

// (* RLOC = "X1Y290" *)
gpc006 gpcL1_290 ({pp18[24],pp19[23],pp20[22],pp21[21],pp22[20],pp23[19]},gpcOutL1_290);
wire [2:0] gpcOutL1_291;

// (* RLOC = "X1Y291" *)
gpc006 gpcL1_291 ({pp24[24],pp25[23],pp26[22],pp27[21],pp28[20],pp29[19]},gpcOutL1_291);
wire [2:0] gpcOutL1_292;

// (* RLOC = "X1Y292" *)
gpc006 gpcL1_292 ({pp30[24],pp31[23],pp32[22],pp33[21],pp34[20],pp35[19]},gpcOutL1_292);
wire [2:0] gpcOutL1_293;

// (* RLOC = "X1Y293" *)
gpc006 gpcL1_293 ({pp36[24],pp37[23],pp38[22],pp39[21],pp40[20],pp41[19]},gpcOutL1_293);
wire [2:0] gpcOutL1_294;

// (* RLOC = "X1Y294" *)
gpc006 gpcL1_294 ({pp39[27],pp40[26],pp41[25],pp42[24],pp43[23],pp44[22]},gpcOutL1_294);
wire [2:0] gpcOutL1_295;

// (* RLOC = "X1Y295" *)
gpc006 gpcL1_295 ({pp39[33],pp40[32],pp41[31],pp42[30],pp43[29],pp44[28]},gpcOutL1_295);
wire [2:0] gpcOutL1_296;

// (* RLOC = "X1Y296" *)
gpc006 gpcL1_296 ({pp39[39],pp40[38],pp41[37],pp42[36],pp43[35],pp44[34]},gpcOutL1_296);
wire [2:0] gpcOutL1_297;

// (* RLOC = "X1Y297" *)
gpc006 gpcL1_297 ({pp39[45],pp40[44],pp41[43],pp42[42],pp43[41],pp44[40]},gpcOutL1_297);
wire [2:0] gpcOutL1_298;

// (* RLOC = "X1Y298" *)
gpc006 gpcL1_298 ({pp39[51],pp40[50],pp41[49],pp42[48],pp43[47],pp44[46]},gpcOutL1_298);
wire [2:0] gpcOutL1_299;

// (* RLOC = "X1Y299" *)
gpc006 gpcL1_299 ({pp39[57],pp40[56],pp41[55],pp42[54],pp43[53],pp44[52]},gpcOutL1_299);
wire [2:0] gpcOutL1_300;

// (* RLOC = "X1Y300" *)
gpc006 gpcL1_300 ({pp39[63],pp40[62],pp41[61],pp42[60],pp43[59],pp44[58]},gpcOutL1_300);
wire [2:0] gpcOutL1_301;

// (* RLOC = "X1Y301" *)
gpc006 gpcL1_301 ({pp0[23],pp1[22],pp2[21],pp3[20],pp4[19],pp5[18]},gpcOutL1_301);
wire [2:0] gpcOutL1_302;

// (* RLOC = "X1Y302" *)
gpc006 gpcL1_302 ({pp6[23],pp7[22],pp8[21],pp9[20],pp10[19],pp11[18]},gpcOutL1_302);
wire [2:0] gpcOutL1_303;

// (* RLOC = "X1Y303" *)
gpc006 gpcL1_303 ({pp12[23],pp13[22],pp14[21],pp15[20],pp16[19],pp17[18]},gpcOutL1_303);
wire [2:0] gpcOutL1_304;

// (* RLOC = "X1Y304" *)
gpc006 gpcL1_304 ({pp18[23],pp19[22],pp20[21],pp21[20],pp22[19],pp23[18]},gpcOutL1_304);
wire [2:0] gpcOutL1_305;

// (* RLOC = "X1Y305" *)
gpc006 gpcL1_305 ({pp24[23],pp25[22],pp26[21],pp27[20],pp28[19],pp29[18]},gpcOutL1_305);
wire [2:0] gpcOutL1_306;

// (* RLOC = "X1Y306" *)
gpc006 gpcL1_306 ({pp30[23],pp31[22],pp32[21],pp33[20],pp34[19],pp35[18]},gpcOutL1_306);
wire [2:0] gpcOutL1_307;

// (* RLOC = "X1Y307" *)
gpc006 gpcL1_307 ({pp36[23],pp37[22],pp38[21],pp39[20],pp40[19],pp41[18]},gpcOutL1_307);
wire [2:0] gpcOutL1_308;

// (* RLOC = "X1Y308" *)
gpc006 gpcL1_308 ({pp40[27],pp41[26],pp42[25],pp43[24],pp44[23],pp45[22]},gpcOutL1_308);
wire [2:0] gpcOutL1_309;

// (* RLOC = "X1Y309" *)
gpc006 gpcL1_309 ({pp40[33],pp41[32],pp42[31],pp43[30],pp44[29],pp45[28]},gpcOutL1_309);
wire [2:0] gpcOutL1_310;

// (* RLOC = "X1Y310" *)
gpc006 gpcL1_310 ({pp40[39],pp41[38],pp42[37],pp43[36],pp44[35],pp45[34]},gpcOutL1_310);
wire [2:0] gpcOutL1_311;

// (* RLOC = "X1Y311" *)
gpc006 gpcL1_311 ({pp40[45],pp41[44],pp42[43],pp43[42],pp44[41],pp45[40]},gpcOutL1_311);
wire [2:0] gpcOutL1_312;

// (* RLOC = "X1Y312" *)
gpc006 gpcL1_312 ({pp40[51],pp41[50],pp42[49],pp43[48],pp44[47],pp45[46]},gpcOutL1_312);
wire [2:0] gpcOutL1_313;

// (* RLOC = "X1Y313" *)
gpc006 gpcL1_313 ({pp40[57],pp41[56],pp42[55],pp43[54],pp44[53],pp45[52]},gpcOutL1_313);
wire [2:0] gpcOutL1_314;

// (* RLOC = "X1Y314" *)
gpc006 gpcL1_314 ({pp40[63],pp41[62],pp42[61],pp43[60],pp44[59],pp45[58]},gpcOutL1_314);
wire [2:0] gpcOutL1_315;

// (* RLOC = "X1Y315" *)
gpc006 gpcL1_315 ({pp0[22],pp1[21],pp2[20],pp3[19],pp4[18],pp5[17]},gpcOutL1_315);
wire [2:0] gpcOutL1_316;

// (* RLOC = "X1Y316" *)
gpc006 gpcL1_316 ({pp6[22],pp7[21],pp8[20],pp9[19],pp10[18],pp11[17]},gpcOutL1_316);
wire [2:0] gpcOutL1_317;

// (* RLOC = "X1Y317" *)
gpc006 gpcL1_317 ({pp12[22],pp13[21],pp14[20],pp15[19],pp16[18],pp17[17]},gpcOutL1_317);
wire [2:0] gpcOutL1_318;

// (* RLOC = "X1Y318" *)
gpc006 gpcL1_318 ({pp18[22],pp19[21],pp20[20],pp21[19],pp22[18],pp23[17]},gpcOutL1_318);
wire [2:0] gpcOutL1_319;

// (* RLOC = "X1Y319" *)
gpc006 gpcL1_319 ({pp24[22],pp25[21],pp26[20],pp27[19],pp28[18],pp29[17]},gpcOutL1_319);
wire [2:0] gpcOutL1_320;

// (* RLOC = "X1Y320" *)
gpc006 gpcL1_320 ({pp30[22],pp31[21],pp32[20],pp33[19],pp34[18],pp35[17]},gpcOutL1_320);
wire [2:0] gpcOutL1_321;

// (* RLOC = "X1Y321" *)
gpc006 gpcL1_321 ({pp36[22],pp37[21],pp38[20],pp39[19],pp40[18],pp41[17]},gpcOutL1_321);
wire [2:0] gpcOutL1_322;

// (* RLOC = "X1Y322" *)
gpc006 gpcL1_322 ({pp41[27],pp42[26],pp43[25],pp44[24],pp45[23],pp46[22]},gpcOutL1_322);
wire [2:0] gpcOutL1_323;

// (* RLOC = "X1Y323" *)
gpc006 gpcL1_323 ({pp41[33],pp42[32],pp43[31],pp44[30],pp45[29],pp46[28]},gpcOutL1_323);
wire [2:0] gpcOutL1_324;

// (* RLOC = "X1Y324" *)
gpc006 gpcL1_324 ({pp41[39],pp42[38],pp43[37],pp44[36],pp45[35],pp46[34]},gpcOutL1_324);
wire [2:0] gpcOutL1_325;

// (* RLOC = "X1Y325" *)
gpc006 gpcL1_325 ({pp41[45],pp42[44],pp43[43],pp44[42],pp45[41],pp46[40]},gpcOutL1_325);
wire [2:0] gpcOutL1_326;

// (* RLOC = "X1Y326" *)
gpc006 gpcL1_326 ({pp41[51],pp42[50],pp43[49],pp44[48],pp45[47],pp46[46]},gpcOutL1_326);
wire [2:0] gpcOutL1_327;

// (* RLOC = "X1Y327" *)
gpc006 gpcL1_327 ({pp41[57],pp42[56],pp43[55],pp44[54],pp45[53],pp46[52]},gpcOutL1_327);
wire [2:0] gpcOutL1_328;

// (* RLOC = "X1Y328" *)
gpc006 gpcL1_328 ({pp41[63],pp42[62],pp43[61],pp44[60],pp45[59],pp46[58]},gpcOutL1_328);
wire [2:0] gpcOutL1_329;

// (* RLOC = "X1Y329" *)
gpc006 gpcL1_329 ({pp0[21],pp1[20],pp2[19],pp3[18],pp4[17],pp5[16]},gpcOutL1_329);
wire [2:0] gpcOutL1_330;

// (* RLOC = "X1Y330" *)
gpc006 gpcL1_330 ({pp6[21],pp7[20],pp8[19],pp9[18],pp10[17],pp11[16]},gpcOutL1_330);
wire [2:0] gpcOutL1_331;

// (* RLOC = "X1Y331" *)
gpc006 gpcL1_331 ({pp12[21],pp13[20],pp14[19],pp15[18],pp16[17],pp17[16]},gpcOutL1_331);
wire [2:0] gpcOutL1_332;

// (* RLOC = "X1Y332" *)
gpc006 gpcL1_332 ({pp18[21],pp19[20],pp20[19],pp21[18],pp22[17],pp23[16]},gpcOutL1_332);
wire [2:0] gpcOutL1_333;

// (* RLOC = "X1Y333" *)
gpc006 gpcL1_333 ({pp24[21],pp25[20],pp26[19],pp27[18],pp28[17],pp29[16]},gpcOutL1_333);
wire [2:0] gpcOutL1_334;

// (* RLOC = "X1Y334" *)
gpc006 gpcL1_334 ({pp30[21],pp31[20],pp32[19],pp33[18],pp34[17],pp35[16]},gpcOutL1_334);
wire [2:0] gpcOutL1_335;

// (* RLOC = "X1Y335" *)
gpc006 gpcL1_335 ({pp36[21],pp37[20],pp38[19],pp39[18],pp40[17],pp41[16]},gpcOutL1_335);
wire [2:0] gpcOutL1_336;

// (* RLOC = "X1Y336" *)
gpc006 gpcL1_336 ({pp42[21],pp43[20],pp44[19],pp45[18],pp46[17],pp47[16]},gpcOutL1_336);
wire [2:0] gpcOutL1_337;

// (* RLOC = "X1Y337" *)
gpc006 gpcL1_337 ({pp42[27],pp43[26],pp44[25],pp45[24],pp46[23],pp47[22]},gpcOutL1_337);
wire [2:0] gpcOutL1_338;

// (* RLOC = "X1Y338" *)
gpc006 gpcL1_338 ({pp42[33],pp43[32],pp44[31],pp45[30],pp46[29],pp47[28]},gpcOutL1_338);
wire [2:0] gpcOutL1_339;

// (* RLOC = "X1Y339" *)
gpc006 gpcL1_339 ({pp42[39],pp43[38],pp44[37],pp45[36],pp46[35],pp47[34]},gpcOutL1_339);
wire [2:0] gpcOutL1_340;

// (* RLOC = "X1Y340" *)
gpc006 gpcL1_340 ({pp42[45],pp43[44],pp44[43],pp45[42],pp46[41],pp47[40]},gpcOutL1_340);
wire [2:0] gpcOutL1_341;

// (* RLOC = "X1Y341" *)
gpc006 gpcL1_341 ({pp42[51],pp43[50],pp44[49],pp45[48],pp46[47],pp47[46]},gpcOutL1_341);
wire [2:0] gpcOutL1_342;

// (* RLOC = "X1Y342" *)
gpc006 gpcL1_342 ({pp42[57],pp43[56],pp44[55],pp45[54],pp46[53],pp47[52]},gpcOutL1_342);
wire [2:0] gpcOutL1_343;

// (* RLOC = "X1Y343" *)
gpc006 gpcL1_343 ({pp42[63],pp43[62],pp44[61],pp45[60],pp46[59],pp47[58]},gpcOutL1_343);
wire [2:0] gpcOutL1_344;

// (* RLOC = "X1Y344" *)
gpc006 gpcL1_344 ({pp0[20],pp1[19],pp2[18],pp3[17],pp4[16],pp5[15]},gpcOutL1_344);
wire [2:0] gpcOutL1_345;

// (* RLOC = "X1Y345" *)
gpc006 gpcL1_345 ({pp6[20],pp7[19],pp8[18],pp9[17],pp10[16],pp11[15]},gpcOutL1_345);
wire [2:0] gpcOutL1_346;

// (* RLOC = "X1Y346" *)
gpc006 gpcL1_346 ({pp12[20],pp13[19],pp14[18],pp15[17],pp16[16],pp17[15]},gpcOutL1_346);
wire [2:0] gpcOutL1_347;

// (* RLOC = "X1Y347" *)
gpc006 gpcL1_347 ({pp18[20],pp19[19],pp20[18],pp21[17],pp22[16],pp23[15]},gpcOutL1_347);
wire [2:0] gpcOutL1_348;

// (* RLOC = "X1Y348" *)
gpc006 gpcL1_348 ({pp24[20],pp25[19],pp26[18],pp27[17],pp28[16],pp29[15]},gpcOutL1_348);
wire [2:0] gpcOutL1_349;

// (* RLOC = "X1Y349" *)
gpc006 gpcL1_349 ({pp30[20],pp31[19],pp32[18],pp33[17],pp34[16],pp35[15]},gpcOutL1_349);
wire [2:0] gpcOutL1_350;

// (* RLOC = "X1Y350" *)
gpc006 gpcL1_350 ({pp36[20],pp37[19],pp38[18],pp39[17],pp40[16],pp41[15]},gpcOutL1_350);
wire [2:0] gpcOutL1_351;

// (* RLOC = "X1Y351" *)
gpc006 gpcL1_351 ({pp42[20],pp43[19],pp44[18],pp45[17],pp46[16],pp47[15]},gpcOutL1_351);
wire [2:0] gpcOutL1_352;

// (* RLOC = "X1Y352" *)
gpc006 gpcL1_352 ({pp43[21],pp44[20],pp45[19],pp46[18],pp47[17],pp48[16]},gpcOutL1_352);
wire [2:0] gpcOutL1_353;

// (* RLOC = "X1Y353" *)
gpc006 gpcL1_353 ({pp43[27],pp44[26],pp45[25],pp46[24],pp47[23],pp48[22]},gpcOutL1_353);
wire [2:0] gpcOutL1_354;

// (* RLOC = "X1Y354" *)
gpc006 gpcL1_354 ({pp43[33],pp44[32],pp45[31],pp46[30],pp47[29],pp48[28]},gpcOutL1_354);
wire [2:0] gpcOutL1_355;

// (* RLOC = "X1Y355" *)
gpc006 gpcL1_355 ({pp43[39],pp44[38],pp45[37],pp46[36],pp47[35],pp48[34]},gpcOutL1_355);
wire [2:0] gpcOutL1_356;

// (* RLOC = "X1Y356" *)
gpc006 gpcL1_356 ({pp43[45],pp44[44],pp45[43],pp46[42],pp47[41],pp48[40]},gpcOutL1_356);
wire [2:0] gpcOutL1_357;

// (* RLOC = "X1Y357" *)
gpc006 gpcL1_357 ({pp43[51],pp44[50],pp45[49],pp46[48],pp47[47],pp48[46]},gpcOutL1_357);
wire [2:0] gpcOutL1_358;

// (* RLOC = "X1Y358" *)
gpc006 gpcL1_358 ({pp43[57],pp44[56],pp45[55],pp46[54],pp47[53],pp48[52]},gpcOutL1_358);
wire [2:0] gpcOutL1_359;

// (* RLOC = "X1Y359" *)
gpc006 gpcL1_359 ({pp43[63],pp44[62],pp45[61],pp46[60],pp47[59],pp48[58]},gpcOutL1_359);
wire [2:0] gpcOutL1_360;

// (* RLOC = "X1Y360" *)
gpc006 gpcL1_360 ({pp0[19],pp1[18],pp2[17],pp3[16],pp4[15],pp5[14]},gpcOutL1_360);
wire [2:0] gpcOutL1_361;

// (* RLOC = "X1Y361" *)
gpc006 gpcL1_361 ({pp6[19],pp7[18],pp8[17],pp9[16],pp10[15],pp11[14]},gpcOutL1_361);
wire [2:0] gpcOutL1_362;

// (* RLOC = "X1Y362" *)
gpc006 gpcL1_362 ({pp12[19],pp13[18],pp14[17],pp15[16],pp16[15],pp17[14]},gpcOutL1_362);
wire [2:0] gpcOutL1_363;

// (* RLOC = "X1Y363" *)
gpc006 gpcL1_363 ({pp18[19],pp19[18],pp20[17],pp21[16],pp22[15],pp23[14]},gpcOutL1_363);
wire [2:0] gpcOutL1_364;

// (* RLOC = "X1Y364" *)
gpc006 gpcL1_364 ({pp24[19],pp25[18],pp26[17],pp27[16],pp28[15],pp29[14]},gpcOutL1_364);
wire [2:0] gpcOutL1_365;

// (* RLOC = "X1Y365" *)
gpc006 gpcL1_365 ({pp30[19],pp31[18],pp32[17],pp33[16],pp34[15],pp35[14]},gpcOutL1_365);
wire [2:0] gpcOutL1_366;

// (* RLOC = "X1Y366" *)
gpc006 gpcL1_366 ({pp36[19],pp37[18],pp38[17],pp39[16],pp40[15],pp41[14]},gpcOutL1_366);
wire [2:0] gpcOutL1_367;

// (* RLOC = "X1Y367" *)
gpc006 gpcL1_367 ({pp42[19],pp43[18],pp44[17],pp45[16],pp46[15],pp47[14]},gpcOutL1_367);
wire [2:0] gpcOutL1_368;

// (* RLOC = "X1Y368" *)
gpc006 gpcL1_368 ({pp44[21],pp45[20],pp46[19],pp47[18],pp48[17],pp49[16]},gpcOutL1_368);
wire [2:0] gpcOutL1_369;

// (* RLOC = "X1Y369" *)
gpc006 gpcL1_369 ({pp44[27],pp45[26],pp46[25],pp47[24],pp48[23],pp49[22]},gpcOutL1_369);
wire [2:0] gpcOutL1_370;

// (* RLOC = "X1Y370" *)
gpc006 gpcL1_370 ({pp44[33],pp45[32],pp46[31],pp47[30],pp48[29],pp49[28]},gpcOutL1_370);
wire [2:0] gpcOutL1_371;

// (* RLOC = "X1Y371" *)
gpc006 gpcL1_371 ({pp44[39],pp45[38],pp46[37],pp47[36],pp48[35],pp49[34]},gpcOutL1_371);
wire [2:0] gpcOutL1_372;

// (* RLOC = "X1Y372" *)
gpc006 gpcL1_372 ({pp44[45],pp45[44],pp46[43],pp47[42],pp48[41],pp49[40]},gpcOutL1_372);
wire [2:0] gpcOutL1_373;

// (* RLOC = "X1Y373" *)
gpc006 gpcL1_373 ({pp44[51],pp45[50],pp46[49],pp47[48],pp48[47],pp49[46]},gpcOutL1_373);
wire [2:0] gpcOutL1_374;

// (* RLOC = "X1Y374" *)
gpc006 gpcL1_374 ({pp44[57],pp45[56],pp46[55],pp47[54],pp48[53],pp49[52]},gpcOutL1_374);
wire [2:0] gpcOutL1_375;

// (* RLOC = "X1Y375" *)
gpc006 gpcL1_375 ({pp44[63],pp45[62],pp46[61],pp47[60],pp48[59],pp49[58]},gpcOutL1_375);
wire [2:0] gpcOutL1_376;

// (* RLOC = "X1Y376" *)
gpc006 gpcL1_376 ({pp0[18],pp1[17],pp2[16],pp3[15],pp4[14],pp5[13]},gpcOutL1_376);
wire [2:0] gpcOutL1_377;

// (* RLOC = "X1Y377" *)
gpc006 gpcL1_377 ({pp6[18],pp7[17],pp8[16],pp9[15],pp10[14],pp11[13]},gpcOutL1_377);
wire [2:0] gpcOutL1_378;

// (* RLOC = "X1Y378" *)
gpc006 gpcL1_378 ({pp12[18],pp13[17],pp14[16],pp15[15],pp16[14],pp17[13]},gpcOutL1_378);
wire [2:0] gpcOutL1_379;

// (* RLOC = "X1Y379" *)
gpc006 gpcL1_379 ({pp18[18],pp19[17],pp20[16],pp21[15],pp22[14],pp23[13]},gpcOutL1_379);
wire [2:0] gpcOutL1_380;

// (* RLOC = "X1Y380" *)
gpc006 gpcL1_380 ({pp24[18],pp25[17],pp26[16],pp27[15],pp28[14],pp29[13]},gpcOutL1_380);
wire [2:0] gpcOutL1_381;

// (* RLOC = "X1Y381" *)
gpc006 gpcL1_381 ({pp30[18],pp31[17],pp32[16],pp33[15],pp34[14],pp35[13]},gpcOutL1_381);
wire [2:0] gpcOutL1_382;

// (* RLOC = "X1Y382" *)
gpc006 gpcL1_382 ({pp36[18],pp37[17],pp38[16],pp39[15],pp40[14],pp41[13]},gpcOutL1_382);
wire [2:0] gpcOutL1_383;

// (* RLOC = "X1Y383" *)
gpc006 gpcL1_383 ({pp42[18],pp43[17],pp44[16],pp45[15],pp46[14],pp47[13]},gpcOutL1_383);
wire [2:0] gpcOutL1_384;

// (* RLOC = "X1Y384" *)
gpc006 gpcL1_384 ({pp45[21],pp46[20],pp47[19],pp48[18],pp49[17],pp50[16]},gpcOutL1_384);
wire [2:0] gpcOutL1_385;

// (* RLOC = "X1Y385" *)
gpc006 gpcL1_385 ({pp45[27],pp46[26],pp47[25],pp48[24],pp49[23],pp50[22]},gpcOutL1_385);
wire [2:0] gpcOutL1_386;

// (* RLOC = "X1Y386" *)
gpc006 gpcL1_386 ({pp45[33],pp46[32],pp47[31],pp48[30],pp49[29],pp50[28]},gpcOutL1_386);
wire [2:0] gpcOutL1_387;

// (* RLOC = "X1Y387" *)
gpc006 gpcL1_387 ({pp45[39],pp46[38],pp47[37],pp48[36],pp49[35],pp50[34]},gpcOutL1_387);
wire [2:0] gpcOutL1_388;

// (* RLOC = "X1Y388" *)
gpc006 gpcL1_388 ({pp45[45],pp46[44],pp47[43],pp48[42],pp49[41],pp50[40]},gpcOutL1_388);
wire [2:0] gpcOutL1_389;

// (* RLOC = "X1Y389" *)
gpc006 gpcL1_389 ({pp45[51],pp46[50],pp47[49],pp48[48],pp49[47],pp50[46]},gpcOutL1_389);
wire [2:0] gpcOutL1_390;

// (* RLOC = "X1Y390" *)
gpc006 gpcL1_390 ({pp45[57],pp46[56],pp47[55],pp48[54],pp49[53],pp50[52]},gpcOutL1_390);
wire [2:0] gpcOutL1_391;

// (* RLOC = "X1Y391" *)
gpc006 gpcL1_391 ({pp45[63],pp46[62],pp47[61],pp48[60],pp49[59],pp50[58]},gpcOutL1_391);
wire [2:0] gpcOutL1_392;

// (* RLOC = "X1Y392" *)
gpc006 gpcL1_392 ({pp0[17],pp1[16],pp2[15],pp3[14],pp4[13],pp5[12]},gpcOutL1_392);
wire [2:0] gpcOutL1_393;

// (* RLOC = "X1Y393" *)
gpc006 gpcL1_393 ({pp6[17],pp7[16],pp8[15],pp9[14],pp10[13],pp11[12]},gpcOutL1_393);
wire [2:0] gpcOutL1_394;

// (* RLOC = "X1Y394" *)
gpc006 gpcL1_394 ({pp12[17],pp13[16],pp14[15],pp15[14],pp16[13],pp17[12]},gpcOutL1_394);
wire [2:0] gpcOutL1_395;

// (* RLOC = "X1Y395" *)
gpc006 gpcL1_395 ({pp18[17],pp19[16],pp20[15],pp21[14],pp22[13],pp23[12]},gpcOutL1_395);
wire [2:0] gpcOutL1_396;

// (* RLOC = "X1Y396" *)
gpc006 gpcL1_396 ({pp24[17],pp25[16],pp26[15],pp27[14],pp28[13],pp29[12]},gpcOutL1_396);
wire [2:0] gpcOutL1_397;

// (* RLOC = "X1Y397" *)
gpc006 gpcL1_397 ({pp30[17],pp31[16],pp32[15],pp33[14],pp34[13],pp35[12]},gpcOutL1_397);
wire [2:0] gpcOutL1_398;

// (* RLOC = "X1Y398" *)
gpc006 gpcL1_398 ({pp36[17],pp37[16],pp38[15],pp39[14],pp40[13],pp41[12]},gpcOutL1_398);
wire [2:0] gpcOutL1_399;

// (* RLOC = "X1Y399" *)
gpc006 gpcL1_399 ({pp42[17],pp43[16],pp44[15],pp45[14],pp46[13],pp47[12]},gpcOutL1_399);
wire [2:0] gpcOutL1_400;

// (* RLOC = "X1Y400" *)
gpc006 gpcL1_400 ({pp46[21],pp47[20],pp48[19],pp49[18],pp50[17],pp51[16]},gpcOutL1_400);
wire [2:0] gpcOutL1_401;

// (* RLOC = "X1Y401" *)
gpc006 gpcL1_401 ({pp46[27],pp47[26],pp48[25],pp49[24],pp50[23],pp51[22]},gpcOutL1_401);
wire [2:0] gpcOutL1_402;

// (* RLOC = "X1Y402" *)
gpc006 gpcL1_402 ({pp46[33],pp47[32],pp48[31],pp49[30],pp50[29],pp51[28]},gpcOutL1_402);
wire [2:0] gpcOutL1_403;

// (* RLOC = "X1Y403" *)
gpc006 gpcL1_403 ({pp46[39],pp47[38],pp48[37],pp49[36],pp50[35],pp51[34]},gpcOutL1_403);
wire [2:0] gpcOutL1_404;

// (* RLOC = "X1Y404" *)
gpc006 gpcL1_404 ({pp46[45],pp47[44],pp48[43],pp49[42],pp50[41],pp51[40]},gpcOutL1_404);
wire [2:0] gpcOutL1_405;

// (* RLOC = "X1Y405" *)
gpc006 gpcL1_405 ({pp46[51],pp47[50],pp48[49],pp49[48],pp50[47],pp51[46]},gpcOutL1_405);
wire [2:0] gpcOutL1_406;

// (* RLOC = "X1Y406" *)
gpc006 gpcL1_406 ({pp46[57],pp47[56],pp48[55],pp49[54],pp50[53],pp51[52]},gpcOutL1_406);
wire [2:0] gpcOutL1_407;

// (* RLOC = "X1Y407" *)
gpc006 gpcL1_407 ({pp46[63],pp47[62],pp48[61],pp49[60],pp50[59],pp51[58]},gpcOutL1_407);
wire [2:0] gpcOutL1_408;

// (* RLOC = "X1Y408" *)
gpc006 gpcL1_408 ({pp0[16],pp1[15],pp2[14],pp3[13],pp4[12],pp5[11]},gpcOutL1_408);
wire [2:0] gpcOutL1_409;

// (* RLOC = "X1Y409" *)
gpc006 gpcL1_409 ({pp6[16],pp7[15],pp8[14],pp9[13],pp10[12],pp11[11]},gpcOutL1_409);
wire [2:0] gpcOutL1_410;

// (* RLOC = "X1Y410" *)
gpc006 gpcL1_410 ({pp12[16],pp13[15],pp14[14],pp15[13],pp16[12],pp17[11]},gpcOutL1_410);
wire [2:0] gpcOutL1_411;

// (* RLOC = "X1Y411" *)
gpc006 gpcL1_411 ({pp18[16],pp19[15],pp20[14],pp21[13],pp22[12],pp23[11]},gpcOutL1_411);
wire [2:0] gpcOutL1_412;

// (* RLOC = "X1Y412" *)
gpc006 gpcL1_412 ({pp24[16],pp25[15],pp26[14],pp27[13],pp28[12],pp29[11]},gpcOutL1_412);
wire [2:0] gpcOutL1_413;

// (* RLOC = "X1Y413" *)
gpc006 gpcL1_413 ({pp30[16],pp31[15],pp32[14],pp33[13],pp34[12],pp35[11]},gpcOutL1_413);
wire [2:0] gpcOutL1_414;

// (* RLOC = "X1Y414" *)
gpc006 gpcL1_414 ({pp36[16],pp37[15],pp38[14],pp39[13],pp40[12],pp41[11]},gpcOutL1_414);
wire [2:0] gpcOutL1_415;

// (* RLOC = "X1Y415" *)
gpc006 gpcL1_415 ({pp42[16],pp43[15],pp44[14],pp45[13],pp46[12],pp47[11]},gpcOutL1_415);
wire [2:0] gpcOutL1_416;

// (* RLOC = "X1Y416" *)
gpc006 gpcL1_416 ({pp47[21],pp48[20],pp49[19],pp50[18],pp51[17],pp52[16]},gpcOutL1_416);
wire [2:0] gpcOutL1_417;

// (* RLOC = "X1Y417" *)
gpc006 gpcL1_417 ({pp47[27],pp48[26],pp49[25],pp50[24],pp51[23],pp52[22]},gpcOutL1_417);
wire [2:0] gpcOutL1_418;

// (* RLOC = "X1Y418" *)
gpc006 gpcL1_418 ({pp47[33],pp48[32],pp49[31],pp50[30],pp51[29],pp52[28]},gpcOutL1_418);
wire [2:0] gpcOutL1_419;

// (* RLOC = "X1Y419" *)
gpc006 gpcL1_419 ({pp47[39],pp48[38],pp49[37],pp50[36],pp51[35],pp52[34]},gpcOutL1_419);
wire [2:0] gpcOutL1_420;

// (* RLOC = "X1Y420" *)
gpc006 gpcL1_420 ({pp47[45],pp48[44],pp49[43],pp50[42],pp51[41],pp52[40]},gpcOutL1_420);
wire [2:0] gpcOutL1_421;

// (* RLOC = "X1Y421" *)
gpc006 gpcL1_421 ({pp47[51],pp48[50],pp49[49],pp50[48],pp51[47],pp52[46]},gpcOutL1_421);
wire [2:0] gpcOutL1_422;

// (* RLOC = "X1Y422" *)
gpc006 gpcL1_422 ({pp47[57],pp48[56],pp49[55],pp50[54],pp51[53],pp52[52]},gpcOutL1_422);
wire [2:0] gpcOutL1_423;

// (* RLOC = "X1Y423" *)
gpc006 gpcL1_423 ({pp47[63],pp48[62],pp49[61],pp50[60],pp51[59],pp52[58]},gpcOutL1_423);
wire [2:0] gpcOutL1_424;

// (* RLOC = "X1Y424" *)
gpc006 gpcL1_424 ({pp0[15],pp1[14],pp2[13],pp3[12],pp4[11],pp5[10]},gpcOutL1_424);
wire [2:0] gpcOutL1_425;

// (* RLOC = "X1Y425" *)
gpc006 gpcL1_425 ({pp6[15],pp7[14],pp8[13],pp9[12],pp10[11],pp11[10]},gpcOutL1_425);
wire [2:0] gpcOutL1_426;

// (* RLOC = "X1Y426" *)
gpc006 gpcL1_426 ({pp12[15],pp13[14],pp14[13],pp15[12],pp16[11],pp17[10]},gpcOutL1_426);
wire [2:0] gpcOutL1_427;

// (* RLOC = "X1Y427" *)
gpc006 gpcL1_427 ({pp18[15],pp19[14],pp20[13],pp21[12],pp22[11],pp23[10]},gpcOutL1_427);
wire [2:0] gpcOutL1_428;

// (* RLOC = "X1Y428" *)
gpc006 gpcL1_428 ({pp24[15],pp25[14],pp26[13],pp27[12],pp28[11],pp29[10]},gpcOutL1_428);
wire [2:0] gpcOutL1_429;

// (* RLOC = "X1Y429" *)
gpc006 gpcL1_429 ({pp30[15],pp31[14],pp32[13],pp33[12],pp34[11],pp35[10]},gpcOutL1_429);
wire [2:0] gpcOutL1_430;

// (* RLOC = "X1Y430" *)
gpc006 gpcL1_430 ({pp36[15],pp37[14],pp38[13],pp39[12],pp40[11],pp41[10]},gpcOutL1_430);
wire [2:0] gpcOutL1_431;

// (* RLOC = "X1Y431" *)
gpc006 gpcL1_431 ({pp42[15],pp43[14],pp44[13],pp45[12],pp46[11],pp47[10]},gpcOutL1_431);
wire [2:0] gpcOutL1_432;

// (* RLOC = "X1Y432" *)
gpc006 gpcL1_432 ({pp48[15],pp49[14],pp50[13],pp51[12],pp52[11],pp53[10]},gpcOutL1_432);
wire [2:0] gpcOutL1_433;

// (* RLOC = "X1Y433" *)
gpc006 gpcL1_433 ({pp48[21],pp49[20],pp50[19],pp51[18],pp52[17],pp53[16]},gpcOutL1_433);
wire [2:0] gpcOutL1_434;

// (* RLOC = "X1Y434" *)
gpc006 gpcL1_434 ({pp48[27],pp49[26],pp50[25],pp51[24],pp52[23],pp53[22]},gpcOutL1_434);
wire [2:0] gpcOutL1_435;

// (* RLOC = "X1Y435" *)
gpc006 gpcL1_435 ({pp48[33],pp49[32],pp50[31],pp51[30],pp52[29],pp53[28]},gpcOutL1_435);
wire [2:0] gpcOutL1_436;

// (* RLOC = "X1Y436" *)
gpc006 gpcL1_436 ({pp48[39],pp49[38],pp50[37],pp51[36],pp52[35],pp53[34]},gpcOutL1_436);
wire [2:0] gpcOutL1_437;

// (* RLOC = "X1Y437" *)
gpc006 gpcL1_437 ({pp48[45],pp49[44],pp50[43],pp51[42],pp52[41],pp53[40]},gpcOutL1_437);
wire [2:0] gpcOutL1_438;

// (* RLOC = "X1Y438" *)
gpc006 gpcL1_438 ({pp48[51],pp49[50],pp50[49],pp51[48],pp52[47],pp53[46]},gpcOutL1_438);
wire [2:0] gpcOutL1_439;

// (* RLOC = "X1Y439" *)
gpc006 gpcL1_439 ({pp48[57],pp49[56],pp50[55],pp51[54],pp52[53],pp53[52]},gpcOutL1_439);
wire [2:0] gpcOutL1_440;

// (* RLOC = "X1Y440" *)
gpc006 gpcL1_440 ({pp48[63],pp49[62],pp50[61],pp51[60],pp52[59],pp53[58]},gpcOutL1_440);
wire [2:0] gpcOutL1_441;

// (* RLOC = "X1Y441" *)
gpc006 gpcL1_441 ({pp0[14],pp1[13],pp2[12],pp3[11],pp4[10],pp5[9]},gpcOutL1_441);
wire [2:0] gpcOutL1_442;

// (* RLOC = "X1Y442" *)
gpc006 gpcL1_442 ({pp6[14],pp7[13],pp8[12],pp9[11],pp10[10],pp11[9]},gpcOutL1_442);
wire [2:0] gpcOutL1_443;

// (* RLOC = "X1Y443" *)
gpc006 gpcL1_443 ({pp12[14],pp13[13],pp14[12],pp15[11],pp16[10],pp17[9]},gpcOutL1_443);
wire [2:0] gpcOutL1_444;

// (* RLOC = "X1Y444" *)
gpc006 gpcL1_444 ({pp18[14],pp19[13],pp20[12],pp21[11],pp22[10],pp23[9]},gpcOutL1_444);
wire [2:0] gpcOutL1_445;

// (* RLOC = "X1Y445" *)
gpc006 gpcL1_445 ({pp24[14],pp25[13],pp26[12],pp27[11],pp28[10],pp29[9]},gpcOutL1_445);
wire [2:0] gpcOutL1_446;

// (* RLOC = "X1Y446" *)
gpc006 gpcL1_446 ({pp30[14],pp31[13],pp32[12],pp33[11],pp34[10],pp35[9]},gpcOutL1_446);
wire [2:0] gpcOutL1_447;

// (* RLOC = "X1Y447" *)
gpc006 gpcL1_447 ({pp36[14],pp37[13],pp38[12],pp39[11],pp40[10],pp41[9]},gpcOutL1_447);
wire [2:0] gpcOutL1_448;

// (* RLOC = "X1Y448" *)
gpc006 gpcL1_448 ({pp42[14],pp43[13],pp44[12],pp45[11],pp46[10],pp47[9]},gpcOutL1_448);
wire [2:0] gpcOutL1_449;

// (* RLOC = "X1Y449" *)
gpc006 gpcL1_449 ({pp48[14],pp49[13],pp50[12],pp51[11],pp52[10],pp53[9]},gpcOutL1_449);
wire [2:0] gpcOutL1_450;

// (* RLOC = "X1Y450" *)
gpc006 gpcL1_450 ({pp49[15],pp50[14],pp51[13],pp52[12],pp53[11],pp54[10]},gpcOutL1_450);
wire [2:0] gpcOutL1_451;

// (* RLOC = "X1Y451" *)
gpc006 gpcL1_451 ({pp49[21],pp50[20],pp51[19],pp52[18],pp53[17],pp54[16]},gpcOutL1_451);
wire [2:0] gpcOutL1_452;

// (* RLOC = "X1Y452" *)
gpc006 gpcL1_452 ({pp49[27],pp50[26],pp51[25],pp52[24],pp53[23],pp54[22]},gpcOutL1_452);
wire [2:0] gpcOutL1_453;

// (* RLOC = "X1Y453" *)
gpc006 gpcL1_453 ({pp49[33],pp50[32],pp51[31],pp52[30],pp53[29],pp54[28]},gpcOutL1_453);
wire [2:0] gpcOutL1_454;

// (* RLOC = "X1Y454" *)
gpc006 gpcL1_454 ({pp49[39],pp50[38],pp51[37],pp52[36],pp53[35],pp54[34]},gpcOutL1_454);
wire [2:0] gpcOutL1_455;

// (* RLOC = "X1Y455" *)
gpc006 gpcL1_455 ({pp49[45],pp50[44],pp51[43],pp52[42],pp53[41],pp54[40]},gpcOutL1_455);
wire [2:0] gpcOutL1_456;

// (* RLOC = "X1Y456" *)
gpc006 gpcL1_456 ({pp49[51],pp50[50],pp51[49],pp52[48],pp53[47],pp54[46]},gpcOutL1_456);
wire [2:0] gpcOutL1_457;

// (* RLOC = "X1Y457" *)
gpc006 gpcL1_457 ({pp49[57],pp50[56],pp51[55],pp52[54],pp53[53],pp54[52]},gpcOutL1_457);
wire [2:0] gpcOutL1_458;

// (* RLOC = "X1Y458" *)
gpc006 gpcL1_458 ({pp49[63],pp50[62],pp51[61],pp52[60],pp53[59],pp54[58]},gpcOutL1_458);
wire [2:0] gpcOutL1_459;

// (* RLOC = "X1Y459" *)
gpc006 gpcL1_459 ({pp0[13],pp1[12],pp2[11],pp3[10],pp4[9],pp5[8]},gpcOutL1_459);
wire [2:0] gpcOutL1_460;

// (* RLOC = "X1Y460" *)
gpc006 gpcL1_460 ({pp6[13],pp7[12],pp8[11],pp9[10],pp10[9],pp11[8]},gpcOutL1_460);
wire [2:0] gpcOutL1_461;

// (* RLOC = "X1Y461" *)
gpc006 gpcL1_461 ({pp12[13],pp13[12],pp14[11],pp15[10],pp16[9],pp17[8]},gpcOutL1_461);
wire [2:0] gpcOutL1_462;

// (* RLOC = "X1Y462" *)
gpc006 gpcL1_462 ({pp18[13],pp19[12],pp20[11],pp21[10],pp22[9],pp23[8]},gpcOutL1_462);
wire [2:0] gpcOutL1_463;

// (* RLOC = "X1Y463" *)
gpc006 gpcL1_463 ({pp24[13],pp25[12],pp26[11],pp27[10],pp28[9],pp29[8]},gpcOutL1_463);
wire [2:0] gpcOutL1_464;

// (* RLOC = "X1Y464" *)
gpc006 gpcL1_464 ({pp30[13],pp31[12],pp32[11],pp33[10],pp34[9],pp35[8]},gpcOutL1_464);
wire [2:0] gpcOutL1_465;

// (* RLOC = "X1Y465" *)
gpc006 gpcL1_465 ({pp36[13],pp37[12],pp38[11],pp39[10],pp40[9],pp41[8]},gpcOutL1_465);
wire [2:0] gpcOutL1_466;

// (* RLOC = "X1Y466" *)
gpc006 gpcL1_466 ({pp42[13],pp43[12],pp44[11],pp45[10],pp46[9],pp47[8]},gpcOutL1_466);
wire [2:0] gpcOutL1_467;

// (* RLOC = "X1Y467" *)
gpc006 gpcL1_467 ({pp48[13],pp49[12],pp50[11],pp51[10],pp52[9],pp53[8]},gpcOutL1_467);
wire [2:0] gpcOutL1_468;

// (* RLOC = "X1Y468" *)
gpc006 gpcL1_468 ({pp50[15],pp51[14],pp52[13],pp53[12],pp54[11],pp55[10]},gpcOutL1_468);
wire [2:0] gpcOutL1_469;

// (* RLOC = "X1Y469" *)
gpc006 gpcL1_469 ({pp50[21],pp51[20],pp52[19],pp53[18],pp54[17],pp55[16]},gpcOutL1_469);
wire [2:0] gpcOutL1_470;

// (* RLOC = "X1Y470" *)
gpc006 gpcL1_470 ({pp50[27],pp51[26],pp52[25],pp53[24],pp54[23],pp55[22]},gpcOutL1_470);
wire [2:0] gpcOutL1_471;

// (* RLOC = "X1Y471" *)
gpc006 gpcL1_471 ({pp50[33],pp51[32],pp52[31],pp53[30],pp54[29],pp55[28]},gpcOutL1_471);
wire [2:0] gpcOutL1_472;

// (* RLOC = "X1Y472" *)
gpc006 gpcL1_472 ({pp50[39],pp51[38],pp52[37],pp53[36],pp54[35],pp55[34]},gpcOutL1_472);
wire [2:0] gpcOutL1_473;

// (* RLOC = "X1Y473" *)
gpc006 gpcL1_473 ({pp50[45],pp51[44],pp52[43],pp53[42],pp54[41],pp55[40]},gpcOutL1_473);
wire [2:0] gpcOutL1_474;

// (* RLOC = "X1Y474" *)
gpc006 gpcL1_474 ({pp50[51],pp51[50],pp52[49],pp53[48],pp54[47],pp55[46]},gpcOutL1_474);
wire [2:0] gpcOutL1_475;

// (* RLOC = "X1Y475" *)
gpc006 gpcL1_475 ({pp50[57],pp51[56],pp52[55],pp53[54],pp54[53],pp55[52]},gpcOutL1_475);
wire [2:0] gpcOutL1_476;

// (* RLOC = "X1Y476" *)
gpc006 gpcL1_476 ({pp50[63],pp51[62],pp52[61],pp53[60],pp54[59],pp55[58]},gpcOutL1_476);
wire [2:0] gpcOutL1_477;

// (* RLOC = "X1Y477" *)
gpc006 gpcL1_477 ({pp0[12],pp1[11],pp2[10],pp3[9],pp4[8],pp5[7]},gpcOutL1_477);
wire [2:0] gpcOutL1_478;

// (* RLOC = "X1Y478" *)
gpc006 gpcL1_478 ({pp6[12],pp7[11],pp8[10],pp9[9],pp10[8],pp11[7]},gpcOutL1_478);
wire [2:0] gpcOutL1_479;

// (* RLOC = "X1Y479" *)
gpc006 gpcL1_479 ({pp12[12],pp13[11],pp14[10],pp15[9],pp16[8],pp17[7]},gpcOutL1_479);
wire [2:0] gpcOutL1_480;

// (* RLOC = "X1Y480" *)
gpc006 gpcL1_480 ({pp18[12],pp19[11],pp20[10],pp21[9],pp22[8],pp23[7]},gpcOutL1_480);
wire [2:0] gpcOutL1_481;

// (* RLOC = "X1Y481" *)
gpc006 gpcL1_481 ({pp24[12],pp25[11],pp26[10],pp27[9],pp28[8],pp29[7]},gpcOutL1_481);
wire [2:0] gpcOutL1_482;

// (* RLOC = "X1Y482" *)
gpc006 gpcL1_482 ({pp30[12],pp31[11],pp32[10],pp33[9],pp34[8],pp35[7]},gpcOutL1_482);
wire [2:0] gpcOutL1_483;

// (* RLOC = "X1Y483" *)
gpc006 gpcL1_483 ({pp36[12],pp37[11],pp38[10],pp39[9],pp40[8],pp41[7]},gpcOutL1_483);
wire [2:0] gpcOutL1_484;

// (* RLOC = "X1Y484" *)
gpc006 gpcL1_484 ({pp42[12],pp43[11],pp44[10],pp45[9],pp46[8],pp47[7]},gpcOutL1_484);
wire [2:0] gpcOutL1_485;

// (* RLOC = "X1Y485" *)
gpc006 gpcL1_485 ({pp48[12],pp49[11],pp50[10],pp51[9],pp52[8],pp53[7]},gpcOutL1_485);
wire [2:0] gpcOutL1_486;

// (* RLOC = "X1Y486" *)
gpc006 gpcL1_486 ({pp51[15],pp52[14],pp53[13],pp54[12],pp55[11],pp56[10]},gpcOutL1_486);
wire [2:0] gpcOutL1_487;

// (* RLOC = "X1Y487" *)
gpc006 gpcL1_487 ({pp51[21],pp52[20],pp53[19],pp54[18],pp55[17],pp56[16]},gpcOutL1_487);
wire [2:0] gpcOutL1_488;

// (* RLOC = "X1Y488" *)
gpc006 gpcL1_488 ({pp51[27],pp52[26],pp53[25],pp54[24],pp55[23],pp56[22]},gpcOutL1_488);
wire [2:0] gpcOutL1_489;

// (* RLOC = "X1Y489" *)
gpc006 gpcL1_489 ({pp51[33],pp52[32],pp53[31],pp54[30],pp55[29],pp56[28]},gpcOutL1_489);
wire [2:0] gpcOutL1_490;

// (* RLOC = "X1Y490" *)
gpc006 gpcL1_490 ({pp51[39],pp52[38],pp53[37],pp54[36],pp55[35],pp56[34]},gpcOutL1_490);
wire [2:0] gpcOutL1_491;

// (* RLOC = "X1Y491" *)
gpc006 gpcL1_491 ({pp51[45],pp52[44],pp53[43],pp54[42],pp55[41],pp56[40]},gpcOutL1_491);
wire [2:0] gpcOutL1_492;

// (* RLOC = "X1Y492" *)
gpc006 gpcL1_492 ({pp51[51],pp52[50],pp53[49],pp54[48],pp55[47],pp56[46]},gpcOutL1_492);
wire [2:0] gpcOutL1_493;

// (* RLOC = "X1Y493" *)
gpc006 gpcL1_493 ({pp51[57],pp52[56],pp53[55],pp54[54],pp55[53],pp56[52]},gpcOutL1_493);
wire [2:0] gpcOutL1_494;

// (* RLOC = "X1Y494" *)
gpc006 gpcL1_494 ({pp51[63],pp52[62],pp53[61],pp54[60],pp55[59],pp56[58]},gpcOutL1_494);
wire [2:0] gpcOutL1_495;

// (* RLOC = "X1Y495" *)
gpc006 gpcL1_495 ({pp0[11],pp1[10],pp2[9],pp3[8],pp4[7],pp5[6]},gpcOutL1_495);
wire [2:0] gpcOutL1_496;

// (* RLOC = "X1Y496" *)
gpc006 gpcL1_496 ({pp6[11],pp7[10],pp8[9],pp9[8],pp10[7],pp11[6]},gpcOutL1_496);
wire [2:0] gpcOutL1_497;

// (* RLOC = "X1Y497" *)
gpc006 gpcL1_497 ({pp12[11],pp13[10],pp14[9],pp15[8],pp16[7],pp17[6]},gpcOutL1_497);
wire [2:0] gpcOutL1_498;

// (* RLOC = "X1Y498" *)
gpc006 gpcL1_498 ({pp18[11],pp19[10],pp20[9],pp21[8],pp22[7],pp23[6]},gpcOutL1_498);
wire [2:0] gpcOutL1_499;

// (* RLOC = "X1Y499" *)
gpc006 gpcL1_499 ({pp24[11],pp25[10],pp26[9],pp27[8],pp28[7],pp29[6]},gpcOutL1_499);
wire [2:0] gpcOutL1_500;

// (* RLOC = "X1Y500" *)
gpc006 gpcL1_500 ({pp30[11],pp31[10],pp32[9],pp33[8],pp34[7],pp35[6]},gpcOutL1_500);
wire [2:0] gpcOutL1_501;

// (* RLOC = "X1Y501" *)
gpc006 gpcL1_501 ({pp36[11],pp37[10],pp38[9],pp39[8],pp40[7],pp41[6]},gpcOutL1_501);
wire [2:0] gpcOutL1_502;

// (* RLOC = "X1Y502" *)
gpc006 gpcL1_502 ({pp42[11],pp43[10],pp44[9],pp45[8],pp46[7],pp47[6]},gpcOutL1_502);
wire [2:0] gpcOutL1_503;

// (* RLOC = "X1Y503" *)
gpc006 gpcL1_503 ({pp48[11],pp49[10],pp50[9],pp51[8],pp52[7],pp53[6]},gpcOutL1_503);
wire [2:0] gpcOutL1_504;

// (* RLOC = "X1Y504" *)
gpc006 gpcL1_504 ({pp52[15],pp53[14],pp54[13],pp55[12],pp56[11],pp57[10]},gpcOutL1_504);
wire [2:0] gpcOutL1_505;

// (* RLOC = "X1Y505" *)
gpc006 gpcL1_505 ({pp52[21],pp53[20],pp54[19],pp55[18],pp56[17],pp57[16]},gpcOutL1_505);
wire [2:0] gpcOutL1_506;

// (* RLOC = "X1Y506" *)
gpc006 gpcL1_506 ({pp52[27],pp53[26],pp54[25],pp55[24],pp56[23],pp57[22]},gpcOutL1_506);
wire [2:0] gpcOutL1_507;

// (* RLOC = "X1Y507" *)
gpc006 gpcL1_507 ({pp52[33],pp53[32],pp54[31],pp55[30],pp56[29],pp57[28]},gpcOutL1_507);
wire [2:0] gpcOutL1_508;

// (* RLOC = "X1Y508" *)
gpc006 gpcL1_508 ({pp52[39],pp53[38],pp54[37],pp55[36],pp56[35],pp57[34]},gpcOutL1_508);
wire [2:0] gpcOutL1_509;

// (* RLOC = "X1Y509" *)
gpc006 gpcL1_509 ({pp52[45],pp53[44],pp54[43],pp55[42],pp56[41],pp57[40]},gpcOutL1_509);
wire [2:0] gpcOutL1_510;

// (* RLOC = "X1Y510" *)
gpc006 gpcL1_510 ({pp52[51],pp53[50],pp54[49],pp55[48],pp56[47],pp57[46]},gpcOutL1_510);
wire [2:0] gpcOutL1_511;

// (* RLOC = "X1Y511" *)
gpc006 gpcL1_511 ({pp52[57],pp53[56],pp54[55],pp55[54],pp56[53],pp57[52]},gpcOutL1_511);
wire [2:0] gpcOutL1_512;

// (* RLOC = "X1Y512" *)
gpc006 gpcL1_512 ({pp52[63],pp53[62],pp54[61],pp55[60],pp56[59],pp57[58]},gpcOutL1_512);
wire [2:0] gpcOutL1_513;

// (* RLOC = "X1Y513" *)
gpc006 gpcL1_513 ({pp0[10],pp1[9],pp2[8],pp3[7],pp4[6],pp5[5]},gpcOutL1_513);
wire [2:0] gpcOutL1_514;

// (* RLOC = "X1Y514" *)
gpc006 gpcL1_514 ({pp6[10],pp7[9],pp8[8],pp9[7],pp10[6],pp11[5]},gpcOutL1_514);
wire [2:0] gpcOutL1_515;

// (* RLOC = "X1Y515" *)
gpc006 gpcL1_515 ({pp12[10],pp13[9],pp14[8],pp15[7],pp16[6],pp17[5]},gpcOutL1_515);
wire [2:0] gpcOutL1_516;

// (* RLOC = "X1Y516" *)
gpc006 gpcL1_516 ({pp18[10],pp19[9],pp20[8],pp21[7],pp22[6],pp23[5]},gpcOutL1_516);
wire [2:0] gpcOutL1_517;

// (* RLOC = "X1Y517" *)
gpc006 gpcL1_517 ({pp24[10],pp25[9],pp26[8],pp27[7],pp28[6],pp29[5]},gpcOutL1_517);
wire [2:0] gpcOutL1_518;

// (* RLOC = "X1Y518" *)
gpc006 gpcL1_518 ({pp30[10],pp31[9],pp32[8],pp33[7],pp34[6],pp35[5]},gpcOutL1_518);
wire [2:0] gpcOutL1_519;

// (* RLOC = "X1Y519" *)
gpc006 gpcL1_519 ({pp36[10],pp37[9],pp38[8],pp39[7],pp40[6],pp41[5]},gpcOutL1_519);
wire [2:0] gpcOutL1_520;

// (* RLOC = "X1Y520" *)
gpc006 gpcL1_520 ({pp42[10],pp43[9],pp44[8],pp45[7],pp46[6],pp47[5]},gpcOutL1_520);
wire [2:0] gpcOutL1_521;

// (* RLOC = "X1Y521" *)
gpc006 gpcL1_521 ({pp48[10],pp49[9],pp50[8],pp51[7],pp52[6],pp53[5]},gpcOutL1_521);
wire [2:0] gpcOutL1_522;

// (* RLOC = "X1Y522" *)
gpc006 gpcL1_522 ({pp53[15],pp54[14],pp55[13],pp56[12],pp57[11],pp58[10]},gpcOutL1_522);
wire [2:0] gpcOutL1_523;

// (* RLOC = "X1Y523" *)
gpc006 gpcL1_523 ({pp53[21],pp54[20],pp55[19],pp56[18],pp57[17],pp58[16]},gpcOutL1_523);
wire [2:0] gpcOutL1_524;

// (* RLOC = "X1Y524" *)
gpc006 gpcL1_524 ({pp53[27],pp54[26],pp55[25],pp56[24],pp57[23],pp58[22]},gpcOutL1_524);
wire [2:0] gpcOutL1_525;

// (* RLOC = "X1Y525" *)
gpc006 gpcL1_525 ({pp53[33],pp54[32],pp55[31],pp56[30],pp57[29],pp58[28]},gpcOutL1_525);
wire [2:0] gpcOutL1_526;

// (* RLOC = "X1Y526" *)
gpc006 gpcL1_526 ({pp53[39],pp54[38],pp55[37],pp56[36],pp57[35],pp58[34]},gpcOutL1_526);
wire [2:0] gpcOutL1_527;

// (* RLOC = "X1Y527" *)
gpc006 gpcL1_527 ({pp53[45],pp54[44],pp55[43],pp56[42],pp57[41],pp58[40]},gpcOutL1_527);
wire [2:0] gpcOutL1_528;

// (* RLOC = "X1Y528" *)
gpc006 gpcL1_528 ({pp53[51],pp54[50],pp55[49],pp56[48],pp57[47],pp58[46]},gpcOutL1_528);
wire [2:0] gpcOutL1_529;

// (* RLOC = "X1Y529" *)
gpc006 gpcL1_529 ({pp53[57],pp54[56],pp55[55],pp56[54],pp57[53],pp58[52]},gpcOutL1_529);
wire [2:0] gpcOutL1_530;

// (* RLOC = "X1Y530" *)
gpc006 gpcL1_530 ({pp53[63],pp54[62],pp55[61],pp56[60],pp57[59],pp58[58]},gpcOutL1_530);
wire [2:0] gpcOutL1_531;

// (* RLOC = "X1Y531" *)
gpc006 gpcL1_531 ({pp0[9],pp1[8],pp2[7],pp3[6],pp4[5],pp5[4]},gpcOutL1_531);
wire [2:0] gpcOutL1_532;

// (* RLOC = "X1Y532" *)
gpc006 gpcL1_532 ({pp6[9],pp7[8],pp8[7],pp9[6],pp10[5],pp11[4]},gpcOutL1_532);
wire [2:0] gpcOutL1_533;

// (* RLOC = "X1Y533" *)
gpc006 gpcL1_533 ({pp12[9],pp13[8],pp14[7],pp15[6],pp16[5],pp17[4]},gpcOutL1_533);
wire [2:0] gpcOutL1_534;

// (* RLOC = "X1Y534" *)
gpc006 gpcL1_534 ({pp18[9],pp19[8],pp20[7],pp21[6],pp22[5],pp23[4]},gpcOutL1_534);
wire [2:0] gpcOutL1_535;

// (* RLOC = "X1Y535" *)
gpc006 gpcL1_535 ({pp24[9],pp25[8],pp26[7],pp27[6],pp28[5],pp29[4]},gpcOutL1_535);
wire [2:0] gpcOutL1_536;

// (* RLOC = "X1Y536" *)
gpc006 gpcL1_536 ({pp30[9],pp31[8],pp32[7],pp33[6],pp34[5],pp35[4]},gpcOutL1_536);
wire [2:0] gpcOutL1_537;

// (* RLOC = "X1Y537" *)
gpc006 gpcL1_537 ({pp36[9],pp37[8],pp38[7],pp39[6],pp40[5],pp41[4]},gpcOutL1_537);
wire [2:0] gpcOutL1_538;

// (* RLOC = "X1Y538" *)
gpc006 gpcL1_538 ({pp42[9],pp43[8],pp44[7],pp45[6],pp46[5],pp47[4]},gpcOutL1_538);
wire [2:0] gpcOutL1_539;

// (* RLOC = "X1Y539" *)
gpc006 gpcL1_539 ({pp48[9],pp49[8],pp50[7],pp51[6],pp52[5],pp53[4]},gpcOutL1_539);
wire [2:0] gpcOutL1_540;

// (* RLOC = "X1Y540" *)
gpc006 gpcL1_540 ({pp54[9],pp55[8],pp56[7],pp57[6],pp58[5],pp59[4]},gpcOutL1_540);
wire [2:0] gpcOutL1_541;

// (* RLOC = "X1Y541" *)
gpc006 gpcL1_541 ({pp54[15],pp55[14],pp56[13],pp57[12],pp58[11],pp59[10]},gpcOutL1_541);
wire [2:0] gpcOutL1_542;

// (* RLOC = "X1Y542" *)
gpc006 gpcL1_542 ({pp54[21],pp55[20],pp56[19],pp57[18],pp58[17],pp59[16]},gpcOutL1_542);
wire [2:0] gpcOutL1_543;

// (* RLOC = "X1Y543" *)
gpc006 gpcL1_543 ({pp54[27],pp55[26],pp56[25],pp57[24],pp58[23],pp59[22]},gpcOutL1_543);
wire [2:0] gpcOutL1_544;

// (* RLOC = "X1Y544" *)
gpc006 gpcL1_544 ({pp54[33],pp55[32],pp56[31],pp57[30],pp58[29],pp59[28]},gpcOutL1_544);
wire [2:0] gpcOutL1_545;

// (* RLOC = "X1Y545" *)
gpc006 gpcL1_545 ({pp54[39],pp55[38],pp56[37],pp57[36],pp58[35],pp59[34]},gpcOutL1_545);
wire [2:0] gpcOutL1_546;

// (* RLOC = "X1Y546" *)
gpc006 gpcL1_546 ({pp54[45],pp55[44],pp56[43],pp57[42],pp58[41],pp59[40]},gpcOutL1_546);
wire [2:0] gpcOutL1_547;

// (* RLOC = "X1Y547" *)
gpc006 gpcL1_547 ({pp54[51],pp55[50],pp56[49],pp57[48],pp58[47],pp59[46]},gpcOutL1_547);
wire [2:0] gpcOutL1_548;

// (* RLOC = "X1Y548" *)
gpc006 gpcL1_548 ({pp54[57],pp55[56],pp56[55],pp57[54],pp58[53],pp59[52]},gpcOutL1_548);
wire [2:0] gpcOutL1_549;

// (* RLOC = "X1Y549" *)
gpc006 gpcL1_549 ({pp54[63],pp55[62],pp56[61],pp57[60],pp58[59],pp59[58]},gpcOutL1_549);
wire [2:0] gpcOutL1_550;

// (* RLOC = "X1Y550" *)
gpc006 gpcL1_550 ({pp0[8],pp1[7],pp2[6],pp3[5],pp4[4],pp5[3]},gpcOutL1_550);
wire [2:0] gpcOutL1_551;

// (* RLOC = "X1Y551" *)
gpc006 gpcL1_551 ({pp6[8],pp7[7],pp8[6],pp9[5],pp10[4],pp11[3]},gpcOutL1_551);
wire [2:0] gpcOutL1_552;

// (* RLOC = "X1Y552" *)
gpc006 gpcL1_552 ({pp12[8],pp13[7],pp14[6],pp15[5],pp16[4],pp17[3]},gpcOutL1_552);
wire [2:0] gpcOutL1_553;

// (* RLOC = "X1Y553" *)
gpc006 gpcL1_553 ({pp18[8],pp19[7],pp20[6],pp21[5],pp22[4],pp23[3]},gpcOutL1_553);
wire [2:0] gpcOutL1_554;

// (* RLOC = "X1Y554" *)
gpc006 gpcL1_554 ({pp24[8],pp25[7],pp26[6],pp27[5],pp28[4],pp29[3]},gpcOutL1_554);
wire [2:0] gpcOutL1_555;

// (* RLOC = "X1Y555" *)
gpc006 gpcL1_555 ({pp30[8],pp31[7],pp32[6],pp33[5],pp34[4],pp35[3]},gpcOutL1_555);
wire [2:0] gpcOutL1_556;

// (* RLOC = "X1Y556" *)
gpc006 gpcL1_556 ({pp36[8],pp37[7],pp38[6],pp39[5],pp40[4],pp41[3]},gpcOutL1_556);
wire [2:0] gpcOutL1_557;

// (* RLOC = "X1Y557" *)
gpc006 gpcL1_557 ({pp42[8],pp43[7],pp44[6],pp45[5],pp46[4],pp47[3]},gpcOutL1_557);
wire [2:0] gpcOutL1_558;

// (* RLOC = "X1Y558" *)
gpc006 gpcL1_558 ({pp48[8],pp49[7],pp50[6],pp51[5],pp52[4],pp53[3]},gpcOutL1_558);
wire [2:0] gpcOutL1_559;

// (* RLOC = "X1Y559" *)
gpc006 gpcL1_559 ({pp54[8],pp55[7],pp56[6],pp57[5],pp58[4],pp59[3]},gpcOutL1_559);
wire [2:0] gpcOutL1_560;

// (* RLOC = "X1Y560" *)
gpc006 gpcL1_560 ({pp55[9],pp56[8],pp57[7],pp58[6],pp59[5],pp60[4]},gpcOutL1_560);
wire [2:0] gpcOutL1_561;

// (* RLOC = "X1Y561" *)
gpc006 gpcL1_561 ({pp55[15],pp56[14],pp57[13],pp58[12],pp59[11],pp60[10]},gpcOutL1_561);
wire [2:0] gpcOutL1_562;

// (* RLOC = "X1Y562" *)
gpc006 gpcL1_562 ({pp55[21],pp56[20],pp57[19],pp58[18],pp59[17],pp60[16]},gpcOutL1_562);
wire [2:0] gpcOutL1_563;

// (* RLOC = "X1Y563" *)
gpc006 gpcL1_563 ({pp55[27],pp56[26],pp57[25],pp58[24],pp59[23],pp60[22]},gpcOutL1_563);
wire [2:0] gpcOutL1_564;

// (* RLOC = "X1Y564" *)
gpc006 gpcL1_564 ({pp55[33],pp56[32],pp57[31],pp58[30],pp59[29],pp60[28]},gpcOutL1_564);
wire [2:0] gpcOutL1_565;

// (* RLOC = "X1Y565" *)
gpc006 gpcL1_565 ({pp55[39],pp56[38],pp57[37],pp58[36],pp59[35],pp60[34]},gpcOutL1_565);
wire [2:0] gpcOutL1_566;

// (* RLOC = "X1Y566" *)
gpc006 gpcL1_566 ({pp55[45],pp56[44],pp57[43],pp58[42],pp59[41],pp60[40]},gpcOutL1_566);
wire [2:0] gpcOutL1_567;

// (* RLOC = "X1Y567" *)
gpc006 gpcL1_567 ({pp55[51],pp56[50],pp57[49],pp58[48],pp59[47],pp60[46]},gpcOutL1_567);
wire [2:0] gpcOutL1_568;

// (* RLOC = "X1Y568" *)
gpc006 gpcL1_568 ({pp55[57],pp56[56],pp57[55],pp58[54],pp59[53],pp60[52]},gpcOutL1_568);
wire [2:0] gpcOutL1_569;

// (* RLOC = "X1Y569" *)
gpc006 gpcL1_569 ({pp55[63],pp56[62],pp57[61],pp58[60],pp59[59],pp60[58]},gpcOutL1_569);
wire [2:0] gpcOutL1_570;

// (* RLOC = "X1Y570" *)
gpc006 gpcL1_570 ({pp0[7],pp1[6],pp2[5],pp3[4],pp4[3],pp5[2]},gpcOutL1_570);
wire [2:0] gpcOutL1_571;

// (* RLOC = "X1Y571" *)
gpc006 gpcL1_571 ({pp6[7],pp7[6],pp8[5],pp9[4],pp10[3],pp11[2]},gpcOutL1_571);
wire [2:0] gpcOutL1_572;

// (* RLOC = "X1Y572" *)
gpc006 gpcL1_572 ({pp12[7],pp13[6],pp14[5],pp15[4],pp16[3],pp17[2]},gpcOutL1_572);
wire [2:0] gpcOutL1_573;

// (* RLOC = "X1Y573" *)
gpc006 gpcL1_573 ({pp18[7],pp19[6],pp20[5],pp21[4],pp22[3],pp23[2]},gpcOutL1_573);
wire [2:0] gpcOutL1_574;

// (* RLOC = "X1Y574" *)
gpc006 gpcL1_574 ({pp24[7],pp25[6],pp26[5],pp27[4],pp28[3],pp29[2]},gpcOutL1_574);
wire [2:0] gpcOutL1_575;

// (* RLOC = "X1Y575" *)
gpc006 gpcL1_575 ({pp30[7],pp31[6],pp32[5],pp33[4],pp34[3],pp35[2]},gpcOutL1_575);
wire [2:0] gpcOutL1_576;

// (* RLOC = "X1Y576" *)
gpc006 gpcL1_576 ({pp36[7],pp37[6],pp38[5],pp39[4],pp40[3],pp41[2]},gpcOutL1_576);
wire [2:0] gpcOutL1_577;

// (* RLOC = "X1Y577" *)
gpc006 gpcL1_577 ({pp42[7],pp43[6],pp44[5],pp45[4],pp46[3],pp47[2]},gpcOutL1_577);
wire [2:0] gpcOutL1_578;

// (* RLOC = "X1Y578" *)
gpc006 gpcL1_578 ({pp48[7],pp49[6],pp50[5],pp51[4],pp52[3],pp53[2]},gpcOutL1_578);
wire [2:0] gpcOutL1_579;

// (* RLOC = "X1Y579" *)
gpc006 gpcL1_579 ({pp54[7],pp55[6],pp56[5],pp57[4],pp58[3],pp59[2]},gpcOutL1_579);
wire [2:0] gpcOutL1_580;

// (* RLOC = "X1Y580" *)
gpc006 gpcL1_580 ({pp56[9],pp57[8],pp58[7],pp59[6],pp60[5],pp61[4]},gpcOutL1_580);
wire [2:0] gpcOutL1_581;

// (* RLOC = "X1Y581" *)
gpc006 gpcL1_581 ({pp56[15],pp57[14],pp58[13],pp59[12],pp60[11],pp61[10]},gpcOutL1_581);
wire [2:0] gpcOutL1_582;

// (* RLOC = "X1Y582" *)
gpc006 gpcL1_582 ({pp56[21],pp57[20],pp58[19],pp59[18],pp60[17],pp61[16]},gpcOutL1_582);
wire [2:0] gpcOutL1_583;

// (* RLOC = "X1Y583" *)
gpc006 gpcL1_583 ({pp56[27],pp57[26],pp58[25],pp59[24],pp60[23],pp61[22]},gpcOutL1_583);
wire [2:0] gpcOutL1_584;

// (* RLOC = "X1Y584" *)
gpc006 gpcL1_584 ({pp56[33],pp57[32],pp58[31],pp59[30],pp60[29],pp61[28]},gpcOutL1_584);
wire [2:0] gpcOutL1_585;

// (* RLOC = "X1Y585" *)
gpc006 gpcL1_585 ({pp56[39],pp57[38],pp58[37],pp59[36],pp60[35],pp61[34]},gpcOutL1_585);
wire [2:0] gpcOutL1_586;

// (* RLOC = "X1Y586" *)
gpc006 gpcL1_586 ({pp56[45],pp57[44],pp58[43],pp59[42],pp60[41],pp61[40]},gpcOutL1_586);
wire [2:0] gpcOutL1_587;

// (* RLOC = "X1Y587" *)
gpc006 gpcL1_587 ({pp56[51],pp57[50],pp58[49],pp59[48],pp60[47],pp61[46]},gpcOutL1_587);
wire [2:0] gpcOutL1_588;

// (* RLOC = "X1Y588" *)
gpc006 gpcL1_588 ({pp56[57],pp57[56],pp58[55],pp59[54],pp60[53],pp61[52]},gpcOutL1_588);
wire [2:0] gpcOutL1_589;

// (* RLOC = "X1Y589" *)
gpc006 gpcL1_589 ({pp56[63],pp57[62],pp58[61],pp59[60],pp60[59],pp61[58]},gpcOutL1_589);
wire [2:0] gpcOutL1_590;

// (* RLOC = "X1Y590" *)
gpc006 gpcL1_590 ({pp0[6],pp1[5],pp2[4],pp3[3],pp4[2],pp5[1]},gpcOutL1_590);
wire [2:0] gpcOutL1_591;

// (* RLOC = "X1Y591" *)
gpc006 gpcL1_591 ({pp6[6],pp7[5],pp8[4],pp9[3],pp10[2],pp11[1]},gpcOutL1_591);
wire [2:0] gpcOutL1_592;

// (* RLOC = "X1Y592" *)
gpc006 gpcL1_592 ({pp12[6],pp13[5],pp14[4],pp15[3],pp16[2],pp17[1]},gpcOutL1_592);
wire [2:0] gpcOutL1_593;

// (* RLOC = "X1Y593" *)
gpc006 gpcL1_593 ({pp18[6],pp19[5],pp20[4],pp21[3],pp22[2],pp23[1]},gpcOutL1_593);
wire [2:0] gpcOutL1_594;

// (* RLOC = "X1Y594" *)
gpc006 gpcL1_594 ({pp24[6],pp25[5],pp26[4],pp27[3],pp28[2],pp29[1]},gpcOutL1_594);
wire [2:0] gpcOutL1_595;

// (* RLOC = "X1Y595" *)
gpc006 gpcL1_595 ({pp30[6],pp31[5],pp32[4],pp33[3],pp34[2],pp35[1]},gpcOutL1_595);
wire [2:0] gpcOutL1_596;

// (* RLOC = "X1Y596" *)
gpc006 gpcL1_596 ({pp36[6],pp37[5],pp38[4],pp39[3],pp40[2],pp41[1]},gpcOutL1_596);
wire [2:0] gpcOutL1_597;

// (* RLOC = "X1Y597" *)
gpc006 gpcL1_597 ({pp42[6],pp43[5],pp44[4],pp45[3],pp46[2],pp47[1]},gpcOutL1_597);
wire [2:0] gpcOutL1_598;

// (* RLOC = "X1Y598" *)
gpc006 gpcL1_598 ({pp48[6],pp49[5],pp50[4],pp51[3],pp52[2],pp53[1]},gpcOutL1_598);
wire [2:0] gpcOutL1_599;

// (* RLOC = "X1Y599" *)
gpc006 gpcL1_599 ({pp54[6],pp55[5],pp56[4],pp57[3],pp58[2],pp59[1]},gpcOutL1_599);
wire [2:0] gpcOutL1_600;

// (* RLOC = "X1Y600" *)
gpc006 gpcL1_600 ({pp57[9],pp58[8],pp59[7],pp60[6],pp61[5],pp62[4]},gpcOutL1_600);
wire [2:0] gpcOutL1_601;

// (* RLOC = "X1Y601" *)
gpc006 gpcL1_601 ({pp57[15],pp58[14],pp59[13],pp60[12],pp61[11],pp62[10]},gpcOutL1_601);
wire [2:0] gpcOutL1_602;

// (* RLOC = "X1Y602" *)
gpc006 gpcL1_602 ({pp57[21],pp58[20],pp59[19],pp60[18],pp61[17],pp62[16]},gpcOutL1_602);
wire [2:0] gpcOutL1_603;

// (* RLOC = "X1Y603" *)
gpc006 gpcL1_603 ({pp57[27],pp58[26],pp59[25],pp60[24],pp61[23],pp62[22]},gpcOutL1_603);
wire [2:0] gpcOutL1_604;

// (* RLOC = "X1Y604" *)
gpc006 gpcL1_604 ({pp57[33],pp58[32],pp59[31],pp60[30],pp61[29],pp62[28]},gpcOutL1_604);
wire [2:0] gpcOutL1_605;

// (* RLOC = "X1Y605" *)
gpc006 gpcL1_605 ({pp57[39],pp58[38],pp59[37],pp60[36],pp61[35],pp62[34]},gpcOutL1_605);
wire [2:0] gpcOutL1_606;

// (* RLOC = "X1Y606" *)
gpc006 gpcL1_606 ({pp57[45],pp58[44],pp59[43],pp60[42],pp61[41],pp62[40]},gpcOutL1_606);
wire [2:0] gpcOutL1_607;

// (* RLOC = "X1Y607" *)
gpc006 gpcL1_607 ({pp57[51],pp58[50],pp59[49],pp60[48],pp61[47],pp62[46]},gpcOutL1_607);
wire [2:0] gpcOutL1_608;

// (* RLOC = "X1Y608" *)
gpc006 gpcL1_608 ({pp57[57],pp58[56],pp59[55],pp60[54],pp61[53],pp62[52]},gpcOutL1_608);
wire [2:0] gpcOutL1_609;

// (* RLOC = "X1Y609" *)
gpc006 gpcL1_609 ({pp57[63],pp58[62],pp59[61],pp60[60],pp61[59],pp62[58]},gpcOutL1_609);
wire [2:0] gpcOutL1_610;

// (* RLOC = "X1Y610" *)
gpc006 gpcL1_610 ({pp0[5],pp1[4],pp2[3],pp3[2],pp4[1],pp5[0]},gpcOutL1_610);
wire [2:0] gpcOutL1_611;

// (* RLOC = "X1Y611" *)
gpc006 gpcL1_611 ({pp6[5],pp7[4],pp8[3],pp9[2],pp10[1],pp11[0]},gpcOutL1_611);
wire [2:0] gpcOutL1_612;

// (* RLOC = "X1Y612" *)
gpc006 gpcL1_612 ({pp12[5],pp13[4],pp14[3],pp15[2],pp16[1],pp17[0]},gpcOutL1_612);
wire [2:0] gpcOutL1_613;

// (* RLOC = "X1Y613" *)
gpc006 gpcL1_613 ({pp18[5],pp19[4],pp20[3],pp21[2],pp22[1],pp23[0]},gpcOutL1_613);
wire [2:0] gpcOutL1_614;

// (* RLOC = "X1Y614" *)
gpc006 gpcL1_614 ({pp24[5],pp25[4],pp26[3],pp27[2],pp28[1],pp29[0]},gpcOutL1_614);
wire [2:0] gpcOutL1_615;

// (* RLOC = "X1Y615" *)
gpc006 gpcL1_615 ({pp30[5],pp31[4],pp32[3],pp33[2],pp34[1],pp35[0]},gpcOutL1_615);
wire [2:0] gpcOutL1_616;

// (* RLOC = "X1Y616" *)
gpc006 gpcL1_616 ({pp36[5],pp37[4],pp38[3],pp39[2],pp40[1],pp41[0]},gpcOutL1_616);
wire [2:0] gpcOutL1_617;

// (* RLOC = "X1Y617" *)
gpc006 gpcL1_617 ({pp42[5],pp43[4],pp44[3],pp45[2],pp46[1],pp47[0]},gpcOutL1_617);
wire [2:0] gpcOutL1_618;

// (* RLOC = "X1Y618" *)
gpc006 gpcL1_618 ({pp48[5],pp49[4],pp50[3],pp51[2],pp52[1],pp53[0]},gpcOutL1_618);
wire [2:0] gpcOutL1_619;

// (* RLOC = "X1Y619" *)
gpc006 gpcL1_619 ({pp54[5],pp55[4],pp56[3],pp57[2],pp58[1],pp59[0]},gpcOutL1_619);
wire [2:0] gpcOutL1_620;

// (* RLOC = "X1Y620" *)
gpc006 gpcL1_620 ({pp58[9],pp59[8],pp60[7],pp61[6],pp62[5],pp63[4]},gpcOutL1_620);
wire [2:0] gpcOutL1_621;

// (* RLOC = "X1Y621" *)
gpc006 gpcL1_621 ({pp58[15],pp59[14],pp60[13],pp61[12],pp62[11],pp63[10]},gpcOutL1_621);
wire [2:0] gpcOutL1_622;

// (* RLOC = "X1Y622" *)
gpc006 gpcL1_622 ({pp58[21],pp59[20],pp60[19],pp61[18],pp62[17],pp63[16]},gpcOutL1_622);
wire [2:0] gpcOutL1_623;

// (* RLOC = "X1Y623" *)
gpc006 gpcL1_623 ({pp58[27],pp59[26],pp60[25],pp61[24],pp62[23],pp63[22]},gpcOutL1_623);
wire [2:0] gpcOutL1_624;

// (* RLOC = "X1Y624" *)
gpc006 gpcL1_624 ({pp58[33],pp59[32],pp60[31],pp61[30],pp62[29],pp63[28]},gpcOutL1_624);
wire [2:0] gpcOutL1_625;

// (* RLOC = "X1Y625" *)
gpc006 gpcL1_625 ({pp58[39],pp59[38],pp60[37],pp61[36],pp62[35],pp63[34]},gpcOutL1_625);
wire [2:0] gpcOutL1_626;

// (* RLOC = "X1Y626" *)
gpc006 gpcL1_626 ({pp58[45],pp59[44],pp60[43],pp61[42],pp62[41],pp63[40]},gpcOutL1_626);
wire [2:0] gpcOutL1_627;

// (* RLOC = "X1Y627" *)
gpc006 gpcL1_627 ({pp58[51],pp59[50],pp60[49],pp61[48],pp62[47],pp63[46]},gpcOutL1_627);
wire [2:0] gpcOutL1_628;

// (* RLOC = "X1Y628" *)
gpc006 gpcL1_628 ({pp58[57],pp59[56],pp60[55],pp61[54],pp62[53],pp63[52]},gpcOutL1_628);
wire [2:0] gpcOutL1_629;

// (* RLOC = "X1Y629" *)
gpc006 gpcL1_629 ({pp58[63],pp59[62],pp60[61],pp61[60],pp62[59],pp63[58]},gpcOutL1_629);
wire [2:0] gpcOutL1_630;

// (* RLOC = "X1Y630" *)
gpc005 gpcL1_630 ({pp0[4],pp1[3],pp2[2],pp3[1],pp4[0]},gpcOutL1_630);
wire [2:0] gpcOutL1_631;

// (* RLOC = "X1Y631" *)
gpc005 gpcL1_631 ({pp6[4],pp7[3],pp8[2],pp9[1],pp10[0]},gpcOutL1_631);
wire [2:0] gpcOutL1_632;

// (* RLOC = "X1Y632" *)
gpc005 gpcL1_632 ({pp12[4],pp13[3],pp14[2],pp15[1],pp16[0]},gpcOutL1_632);
wire [2:0] gpcOutL1_633;

// (* RLOC = "X1Y633" *)
gpc005 gpcL1_633 ({pp18[4],pp19[3],pp20[2],pp21[1],pp22[0]},gpcOutL1_633);
wire [2:0] gpcOutL1_634;

// (* RLOC = "X1Y634" *)
gpc005 gpcL1_634 ({pp24[4],pp25[3],pp26[2],pp27[1],pp28[0]},gpcOutL1_634);
wire [2:0] gpcOutL1_635;

// (* RLOC = "X1Y635" *)
gpc005 gpcL1_635 ({pp30[4],pp31[3],pp32[2],pp33[1],pp34[0]},gpcOutL1_635);
wire [2:0] gpcOutL1_636;

// (* RLOC = "X1Y636" *)
gpc005 gpcL1_636 ({pp36[4],pp37[3],pp38[2],pp39[1],pp40[0]},gpcOutL1_636);
wire [2:0] gpcOutL1_637;

// (* RLOC = "X1Y637" *)
gpc005 gpcL1_637 ({pp42[4],pp43[3],pp44[2],pp45[1],pp46[0]},gpcOutL1_637);
wire [2:0] gpcOutL1_638;

// (* RLOC = "X1Y638" *)
gpc005 gpcL1_638 ({pp48[4],pp49[3],pp50[2],pp51[1],pp52[0]},gpcOutL1_638);
wire [2:0] gpcOutL1_639;

// (* RLOC = "X1Y639" *)
gpc005 gpcL1_639 ({pp54[4],pp55[3],pp56[2],pp57[1],pp58[0]},gpcOutL1_639);
wire [2:0] gpcOutL1_640;

// (* RLOC = "X1Y640" *)
gpc015 gpcL1_640 ({pp60[9],pp59[9],pp60[8],pp61[7],pp62[6],pp63[5]},gpcOutL1_640);
wire [2:0] gpcOutL1_641;

// (* RLOC = "X1Y641" *)
gpc015 gpcL1_641 ({pp60[15],pp59[15],pp60[14],pp61[13],pp62[12],pp63[11]},gpcOutL1_641);
wire [2:0] gpcOutL1_642;

// (* RLOC = "X1Y642" *)
gpc015 gpcL1_642 ({pp60[21],pp59[21],pp60[20],pp61[19],pp62[18],pp63[17]},gpcOutL1_642);
wire [2:0] gpcOutL1_643;

// (* RLOC = "X1Y643" *)
gpc015 gpcL1_643 ({pp60[27],pp59[27],pp60[26],pp61[25],pp62[24],pp63[23]},gpcOutL1_643);
wire [2:0] gpcOutL1_644;

// (* RLOC = "X1Y644" *)
gpc015 gpcL1_644 ({pp60[33],pp59[33],pp60[32],pp61[31],pp62[30],pp63[29]},gpcOutL1_644);
wire [2:0] gpcOutL1_645;

// (* RLOC = "X1Y645" *)
gpc015 gpcL1_645 ({pp60[39],pp59[39],pp60[38],pp61[37],pp62[36],pp63[35]},gpcOutL1_645);
wire [2:0] gpcOutL1_646;

// (* RLOC = "X1Y646" *)
gpc015 gpcL1_646 ({pp60[45],pp59[45],pp60[44],pp61[43],pp62[42],pp63[41]},gpcOutL1_646);
wire [2:0] gpcOutL1_647;

// (* RLOC = "X1Y647" *)
gpc015 gpcL1_647 ({pp60[51],pp59[51],pp60[50],pp61[49],pp62[48],pp63[47]},gpcOutL1_647);
wire [2:0] gpcOutL1_648;

// (* RLOC = "X1Y648" *)
gpc015 gpcL1_648 ({pp60[57],pp59[57],pp60[56],pp61[55],pp62[54],pp63[53]},gpcOutL1_648);
wire [2:0] gpcOutL1_649;

// (* RLOC = "X1Y649" *)
gpc015 gpcL1_649 ({pp60[63],pp59[63],pp60[62],pp61[61],pp62[60],pp63[59]},gpcOutL1_649);
wire [2:0] gpcOutL1_650;

// (* RLOC = "X1Y650" *)
gpc023 gpcL1_650 ({pp0[3],pp1[2],pp0[2],pp1[1],pp2[0]},gpcOutL1_650);
wire [2:0] gpcOutL1_651;

// (* RLOC = "X1Y651" *)
gpc023 gpcL1_651 ({pp6[3],pp7[2],pp6[2],pp7[1],pp8[0]},gpcOutL1_651);
wire [2:0] gpcOutL1_652;

// (* RLOC = "X1Y652" *)
gpc023 gpcL1_652 ({pp12[3],pp13[2],pp12[2],pp13[1],pp14[0]},gpcOutL1_652);
wire [2:0] gpcOutL1_653;

// (* RLOC = "X1Y653" *)
gpc023 gpcL1_653 ({pp18[3],pp19[2],pp18[2],pp19[1],pp20[0]},gpcOutL1_653);
wire [2:0] gpcOutL1_654;

// (* RLOC = "X1Y654" *)
gpc023 gpcL1_654 ({pp24[3],pp25[2],pp24[2],pp25[1],pp26[0]},gpcOutL1_654);
wire [2:0] gpcOutL1_655;

// (* RLOC = "X1Y655" *)
gpc023 gpcL1_655 ({pp30[3],pp31[2],pp30[2],pp31[1],pp32[0]},gpcOutL1_655);
wire [2:0] gpcOutL1_656;

// (* RLOC = "X1Y656" *)
gpc023 gpcL1_656 ({pp36[3],pp37[2],pp36[2],pp37[1],pp38[0]},gpcOutL1_656);
wire [2:0] gpcOutL1_657;

// (* RLOC = "X1Y657" *)
gpc023 gpcL1_657 ({pp42[3],pp43[2],pp42[2],pp43[1],pp44[0]},gpcOutL1_657);
wire [2:0] gpcOutL1_658;

// (* RLOC = "X1Y658" *)
gpc023 gpcL1_658 ({pp48[3],pp49[2],pp48[2],pp49[1],pp50[0]},gpcOutL1_658);
wire [2:0] gpcOutL1_659;

// (* RLOC = "X1Y659" *)
gpc023 gpcL1_659 ({pp54[3],pp55[2],pp54[2],pp55[1],pp56[0]},gpcOutL1_659);
wire [2:0] gpcOutL1_660;

// (* RLOC = "X1Y660" *)
gpc014 gpcL1_660 ({pp61[3],pp60[3],pp61[2],pp62[1],pp63[0]},gpcOutL1_660);
wire [1:0] gpcOutL1_661;

// (* RLOC = "X1Y661" *)
gpc003 gpcL1_661 ({pp60[2],pp61[1],pp62[0]},gpcOutL1_661);
wire [2:0] gpcOutL1_662;

// (* RLOC = "X1Y662" *)
gpc023 gpcL1_662 ({pp61[9],pp62[8],pp61[8],pp62[7],pp63[6]},gpcOutL1_662);
wire [2:0] gpcOutL1_663;

// (* RLOC = "X1Y663" *)
gpc023 gpcL1_663 ({pp61[15],pp62[14],pp61[14],pp62[13],pp63[12]},gpcOutL1_663);
wire [2:0] gpcOutL1_664;

// (* RLOC = "X1Y664" *)
gpc023 gpcL1_664 ({pp61[21],pp62[20],pp61[20],pp62[19],pp63[18]},gpcOutL1_664);
wire [2:0] gpcOutL1_665;

// (* RLOC = "X1Y665" *)
gpc023 gpcL1_665 ({pp61[27],pp62[26],pp61[26],pp62[25],pp63[24]},gpcOutL1_665);
wire [2:0] gpcOutL1_666;

// (* RLOC = "X1Y666" *)
gpc023 gpcL1_666 ({pp61[33],pp62[32],pp61[32],pp62[31],pp63[30]},gpcOutL1_666);
wire [2:0] gpcOutL1_667;

// (* RLOC = "X1Y667" *)
gpc023 gpcL1_667 ({pp61[39],pp62[38],pp61[38],pp62[37],pp63[36]},gpcOutL1_667);
wire [2:0] gpcOutL1_668;

// (* RLOC = "X1Y668" *)
gpc023 gpcL1_668 ({pp61[45],pp62[44],pp61[44],pp62[43],pp63[42]},gpcOutL1_668);
wire [2:0] gpcOutL1_669;

// (* RLOC = "X1Y669" *)
gpc023 gpcL1_669 ({pp61[51],pp62[50],pp61[50],pp62[49],pp63[48]},gpcOutL1_669);
wire [2:0] gpcOutL1_670;

// (* RLOC = "X1Y670" *)
gpc023 gpcL1_670 ({pp61[57],pp62[56],pp61[56],pp62[55],pp63[54]},gpcOutL1_670);
wire [2:0] gpcOutL1_671;

// (* RLOC = "X1Y671" *)
gpc023 gpcL1_671 ({pp61[63],pp62[62],pp61[62],pp62[61],pp63[60]},gpcOutL1_671);
wire [2:0] gpcOutL1_672;

// (* RLOC = "X1Y672" *)
gpc022 gpcL1_672 ({pp62[3],pp63[2],pp62[2],pp63[1]},gpcOutL1_672);
wire [2:0] gpcOutL2_0;

// (* RLOC = "X2Y0" *)
gpc006 gpcL2_0 ({gpcOutL1_3[0],gpcOutL1_5[1],gpcOutL1_7[2],gpcOutL1_19[0],gpcOutL1_23[1],gpcOutL1_27[2]},gpcOutL2_0);
wire [2:0] gpcOutL2_1;

// (* RLOC = "X2Y1" *)
gpc006 gpcL2_1 ({gpcOutL1_0[0],gpcOutL1_1[1],gpcOutL1_3[2],gpcOutL1_12[0],gpcOutL1_15[1],gpcOutL1_19[2]},gpcOutL2_1);
wire [2:0] gpcOutL2_2;

// (* RLOC = "X2Y2" *)
gpc006 gpcL2_2 ({gpcOutL1_0[1],gpcOutL1_1[2],gpcOutL1_2[0],gpcOutL1_12[1],gpcOutL1_15[2],gpcOutL1_16[0]},gpcOutL2_2);
wire [2:0] gpcOutL2_3;

// (* RLOC = "X2Y3" *)
gpc006 gpcL2_3 ({gpcOutL1_0[2],gpcOutL1_2[1],gpcOutL1_4[0],gpcOutL1_12[2],gpcOutL1_16[1],gpcOutL1_20[0]},gpcOutL2_3);
wire [2:0] gpcOutL2_4;

// (* RLOC = "X2Y4" *)
gpc006 gpcL2_4 ({gpcOutL1_2[2],gpcOutL1_4[1],gpcOutL1_6[0],gpcOutL1_16[2],gpcOutL1_20[1],gpcOutL1_24[0]},gpcOutL2_4);
wire [2:0] gpcOutL2_5;

// (* RLOC = "X2Y5" *)
gpc006 gpcL2_5 ({gpcOutL1_5[0],gpcOutL1_7[1],gpcOutL1_9[2],gpcOutL1_23[0],gpcOutL1_27[1],gpcOutL1_31[2]},gpcOutL2_5);
wire [2:0] gpcOutL2_6;

// (* RLOC = "X2Y6" *)
gpc006 gpcL2_6 ({gpcOutL1_1[0],gpcOutL1_3[1],gpcOutL1_5[2],gpcOutL1_15[0],gpcOutL1_19[1],gpcOutL1_23[2]},gpcOutL2_6);
wire [2:0] gpcOutL2_7;

// (* RLOC = "X2Y7" *)
gpc006 gpcL2_7 ({gpcOutL1_11[0],gpcOutL1_14[1],gpcOutL1_18[2],gpcOutL1_35[0],gpcOutL1_40[1],gpcOutL1_46[2]},gpcOutL2_7);
wire [2:0] gpcOutL2_8;

// (* RLOC = "X2Y8" *)
gpc006 gpcL2_8 ({gpcOutL1_4[2],gpcOutL1_6[1],gpcOutL1_8[0],gpcOutL1_20[2],gpcOutL1_24[1],gpcOutL1_28[0]},gpcOutL2_8);
wire [2:0] gpcOutL2_9;

// (* RLOC = "X2Y9" *)
gpc006 gpcL2_9 ({gpcOutL1_6[2],gpcOutL1_8[1],gpcOutL1_10[0],gpcOutL1_24[2],gpcOutL1_28[1],gpcOutL1_32[0]},gpcOutL2_9);
wire [2:0] gpcOutL2_10;

// (* RLOC = "X2Y10" *)
gpc006 gpcL2_10 ({gpcOutL1_8[2],gpcOutL1_10[1],gpcOutL1_13[0],gpcOutL1_28[2],gpcOutL1_32[1],gpcOutL1_37[0]},gpcOutL2_10);
wire [2:0] gpcOutL2_11;

// (* RLOC = "X2Y11" *)
gpc006 gpcL2_11 ({gpcOutL1_10[2],gpcOutL1_13[1],gpcOutL1_17[0],gpcOutL1_32[2],gpcOutL1_37[1],gpcOutL1_43[0]},gpcOutL2_11);
wire [2:0] gpcOutL2_12;

// (* RLOC = "X2Y12" *)
gpc006 gpcL2_12 ({gpcOutL1_13[2],gpcOutL1_17[1],gpcOutL1_21[0],gpcOutL1_37[2],gpcOutL1_43[1],gpcOutL1_49[0]},gpcOutL2_12);
wire [2:0] gpcOutL2_13;

// (* RLOC = "X2Y13" *)
gpc006 gpcL2_13 ({gpcOutL1_18[0],gpcOutL1_22[1],gpcOutL1_26[2],gpcOutL1_46[0],gpcOutL1_52[1],gpcOutL1_58[2]},gpcOutL2_13);
wire [2:0] gpcOutL2_14;

// (* RLOC = "X2Y14" *)
gpc006 gpcL2_14 ({gpcOutL1_9[0],gpcOutL1_11[1],gpcOutL1_14[2],gpcOutL1_31[0],gpcOutL1_35[1],gpcOutL1_40[2]},gpcOutL2_14);
wire [2:0] gpcOutL2_15;

// (* RLOC = "X2Y15" *)
gpc006 gpcL2_15 ({gpcOutL1_7[0],gpcOutL1_9[1],gpcOutL1_11[2],gpcOutL1_27[0],gpcOutL1_31[1],gpcOutL1_35[2]},gpcOutL2_15);
wire [2:0] gpcOutL2_16;

// (* RLOC = "X2Y16" *)
gpc006 gpcL2_16 ({gpcOutL1_22[0],gpcOutL1_26[1],gpcOutL1_30[2],gpcOutL1_52[0],gpcOutL1_58[1],gpcOutL1_64[2]},gpcOutL2_16);
wire [2:0] gpcOutL2_17;

// (* RLOC = "X2Y17" *)
gpc006 gpcL2_17 ({gpcOutL1_14[0],gpcOutL1_18[1],gpcOutL1_22[2],gpcOutL1_40[0],gpcOutL1_46[1],gpcOutL1_52[2]},gpcOutL2_17);
wire [2:0] gpcOutL2_18;

// (* RLOC = "X2Y18" *)
gpc006 gpcL2_18 ({gpcOutL1_17[2],gpcOutL1_21[1],gpcOutL1_25[0],gpcOutL1_43[2],gpcOutL1_49[1],gpcOutL1_55[0]},gpcOutL2_18);
wire [2:0] gpcOutL2_19;

// (* RLOC = "X2Y19" *)
gpc006 gpcL2_19 ({gpcOutL1_34[0],gpcOutL1_39[1],gpcOutL1_45[2],gpcOutL1_70[0],gpcOutL1_77[1],gpcOutL1_85[2]},gpcOutL2_19);
wire [2:0] gpcOutL2_20;

// (* RLOC = "X2Y20" *)
gpc006 gpcL2_20 ({gpcOutL1_21[2],gpcOutL1_25[1],gpcOutL1_29[0],gpcOutL1_49[2],gpcOutL1_55[1],gpcOutL1_61[0]},gpcOutL2_20);
wire [2:0] gpcOutL2_21;

// (* RLOC = "X2Y21" *)
gpc006 gpcL2_21 ({gpcOutL1_25[2],gpcOutL1_29[1],gpcOutL1_33[0],gpcOutL1_55[2],gpcOutL1_61[1],gpcOutL1_67[0]},gpcOutL2_21);
wire [2:0] gpcOutL2_22;

// (* RLOC = "X2Y22" *)
gpc006 gpcL2_22 ({gpcOutL1_29[2],gpcOutL1_33[1],gpcOutL1_38[0],gpcOutL1_61[2],gpcOutL1_67[1],gpcOutL1_74[0]},gpcOutL2_22);
wire [2:0] gpcOutL2_23;

// (* RLOC = "X2Y23" *)
gpc006 gpcL2_23 ({gpcOutL1_33[2],gpcOutL1_38[1],gpcOutL1_44[0],gpcOutL1_67[2],gpcOutL1_74[1],gpcOutL1_82[0]},gpcOutL2_23);
wire [2:0] gpcOutL2_24;

// (* RLOC = "X2Y24" *)
gpc006 gpcL2_24 ({gpcOutL1_38[2],gpcOutL1_44[1],gpcOutL1_50[0],gpcOutL1_74[2],gpcOutL1_82[1],gpcOutL1_90[0]},gpcOutL2_24);
wire [2:0] gpcOutL2_25;

// (* RLOC = "X2Y25" *)
gpc006 gpcL2_25 ({gpcOutL1_45[0],gpcOutL1_51[1],gpcOutL1_57[2],gpcOutL1_85[0],gpcOutL1_93[1],gpcOutL1_101[2]},gpcOutL2_25);
wire [2:0] gpcOutL2_26;

// (* RLOC = "X2Y26" *)
gpc006 gpcL2_26 ({gpcOutL1_30[0],gpcOutL1_34[1],gpcOutL1_39[2],gpcOutL1_64[0],gpcOutL1_70[1],gpcOutL1_77[2]},gpcOutL2_26);
wire [2:0] gpcOutL2_27;

// (* RLOC = "X2Y27" *)
gpc006 gpcL2_27 ({gpcOutL1_26[0],gpcOutL1_30[1],gpcOutL1_34[2],gpcOutL1_58[0],gpcOutL1_64[1],gpcOutL1_70[2]},gpcOutL2_27);
wire [2:0] gpcOutL2_28;

// (* RLOC = "X2Y28" *)
gpc006 gpcL2_28 ({gpcOutL1_47[0],gpcOutL1_53[1],gpcOutL1_59[2],gpcOutL1_87[0],gpcOutL1_95[1],gpcOutL1_103[2]},gpcOutL2_28);
wire [2:0] gpcOutL2_29;

// (* RLOC = "X2Y29" *)
gpc006 gpcL2_29 ({gpcOutL1_36[0],gpcOutL1_41[1],gpcOutL1_47[2],gpcOutL1_72[0],gpcOutL1_79[1],gpcOutL1_87[2]},gpcOutL2_29);
wire [2:0] gpcOutL2_30;

// (* RLOC = "X2Y30" *)
gpc006 gpcL2_30 ({gpcOutL1_36[1],gpcOutL1_41[2],gpcOutL1_42[0],gpcOutL1_72[1],gpcOutL1_79[2],gpcOutL1_80[0]},gpcOutL2_30);
wire [2:0] gpcOutL2_31;

// (* RLOC = "X2Y31" *)
gpc006 gpcL2_31 ({gpcOutL1_36[2],gpcOutL1_42[1],gpcOutL1_48[0],gpcOutL1_72[2],gpcOutL1_80[1],gpcOutL1_88[0]},gpcOutL2_31);
wire [2:0] gpcOutL2_32;

// (* RLOC = "X2Y32" *)
gpc006 gpcL2_32 ({gpcOutL1_42[2],gpcOutL1_48[1],gpcOutL1_54[0],gpcOutL1_80[2],gpcOutL1_88[1],gpcOutL1_96[0]},gpcOutL2_32);
wire [2:0] gpcOutL2_33;

// (* RLOC = "X2Y33" *)
gpc006 gpcL2_33 ({gpcOutL1_51[0],gpcOutL1_57[1],gpcOutL1_63[2],gpcOutL1_93[0],gpcOutL1_101[1],gpcOutL1_109[2]},gpcOutL2_33);
wire [2:0] gpcOutL2_34;

// (* RLOC = "X2Y34" *)
gpc006 gpcL2_34 ({gpcOutL1_39[0],gpcOutL1_45[1],gpcOutL1_51[2],gpcOutL1_77[0],gpcOutL1_85[1],gpcOutL1_93[2]},gpcOutL2_34);
wire [2:0] gpcOutL2_35;

// (* RLOC = "X2Y35" *)
gpc006 gpcL2_35 ({gpcOutL1_53[0],gpcOutL1_59[1],gpcOutL1_65[2],gpcOutL1_95[0],gpcOutL1_103[1],gpcOutL1_111[2]},gpcOutL2_35);
wire [2:0] gpcOutL2_36;

// (* RLOC = "X2Y36" *)
gpc006 gpcL2_36 ({gpcOutL1_41[0],gpcOutL1_47[1],gpcOutL1_53[2],gpcOutL1_79[0],gpcOutL1_87[1],gpcOutL1_95[2]},gpcOutL2_36);
wire [2:0] gpcOutL2_37;

// (* RLOC = "X2Y37" *)
gpc006 gpcL2_37 ({gpcOutL1_44[2],gpcOutL1_50[1],gpcOutL1_56[0],gpcOutL1_82[2],gpcOutL1_90[1],gpcOutL1_98[0]},gpcOutL2_37);
wire [2:0] gpcOutL2_38;

// (* RLOC = "X2Y38" *)
gpc006 gpcL2_38 ({gpcOutL1_69[0],gpcOutL1_76[1],gpcOutL1_84[2],gpcOutL1_117[0],gpcOutL1_126[1],gpcOutL1_136[2]},gpcOutL2_38);
wire [2:0] gpcOutL2_39;

// (* RLOC = "X2Y39" *)
gpc006 gpcL2_39 ({gpcOutL1_71[0],gpcOutL1_78[1],gpcOutL1_86[2],gpcOutL1_119[0],gpcOutL1_128[1],gpcOutL1_138[2]},gpcOutL2_39);
wire [2:0] gpcOutL2_40;

// (* RLOC = "X2Y40" *)
gpc006 gpcL2_40 ({gpcOutL1_48[2],gpcOutL1_54[1],gpcOutL1_60[0],gpcOutL1_88[2],gpcOutL1_96[1],gpcOutL1_104[0]},gpcOutL2_40);
wire [2:0] gpcOutL2_41;

// (* RLOC = "X2Y41" *)
gpc006 gpcL2_41 ({gpcOutL1_54[2],gpcOutL1_60[1],gpcOutL1_66[0],gpcOutL1_96[2],gpcOutL1_104[1],gpcOutL1_112[0]},gpcOutL2_41);
wire [2:0] gpcOutL2_42;

// (* RLOC = "X2Y42" *)
gpc006 gpcL2_42 ({gpcOutL1_60[2],gpcOutL1_66[1],gpcOutL1_73[0],gpcOutL1_104[2],gpcOutL1_112[1],gpcOutL1_121[0]},gpcOutL2_42);
wire [2:0] gpcOutL2_43;

// (* RLOC = "X2Y43" *)
gpc006 gpcL2_43 ({gpcOutL1_66[2],gpcOutL1_73[1],gpcOutL1_81[0],gpcOutL1_112[2],gpcOutL1_121[1],gpcOutL1_131[0]},gpcOutL2_43);
wire [2:0] gpcOutL2_44;

// (* RLOC = "X2Y44" *)
gpc006 gpcL2_44 ({gpcOutL1_73[2],gpcOutL1_81[1],gpcOutL1_89[0],gpcOutL1_121[2],gpcOutL1_131[1],gpcOutL1_141[0]},gpcOutL2_44);
wire [2:0] gpcOutL2_45;

// (* RLOC = "X2Y45" *)
gpc006 gpcL2_45 ({gpcOutL1_50[2],gpcOutL1_56[1],gpcOutL1_62[0],gpcOutL1_90[2],gpcOutL1_98[1],gpcOutL1_106[0]},gpcOutL2_45);
wire [2:0] gpcOutL2_46;

// (* RLOC = "X2Y46" *)
gpc006 gpcL2_46 ({gpcOutL1_56[2],gpcOutL1_62[1],gpcOutL1_68[0],gpcOutL1_98[2],gpcOutL1_106[1],gpcOutL1_114[0]},gpcOutL2_46);
wire [2:0] gpcOutL2_47;

// (* RLOC = "X2Y47" *)
gpc006 gpcL2_47 ({gpcOutL1_62[2],gpcOutL1_68[1],gpcOutL1_75[0],gpcOutL1_106[2],gpcOutL1_114[1],gpcOutL1_123[0]},gpcOutL2_47);
wire [2:0] gpcOutL2_48;

// (* RLOC = "X2Y48" *)
gpc006 gpcL2_48 ({gpcOutL1_68[2],gpcOutL1_75[1],gpcOutL1_83[0],gpcOutL1_114[2],gpcOutL1_123[1],gpcOutL1_133[0]},gpcOutL2_48);
wire [2:0] gpcOutL2_49;

// (* RLOC = "X2Y49" *)
gpc006 gpcL2_49 ({gpcOutL1_75[2],gpcOutL1_83[1],gpcOutL1_91[0],gpcOutL1_123[2],gpcOutL1_133[1],gpcOutL1_143[0]},gpcOutL2_49);
wire [2:0] gpcOutL2_50;

// (* RLOC = "X2Y50" *)
gpc006 gpcL2_50 ({gpcOutL1_84[0],gpcOutL1_92[1],gpcOutL1_100[2],gpcOutL1_136[0],gpcOutL1_146[1],gpcOutL1_156[2]},gpcOutL2_50);
wire [2:0] gpcOutL2_51;

// (* RLOC = "X2Y51" *)
gpc006 gpcL2_51 ({gpcOutL1_63[0],gpcOutL1_69[1],gpcOutL1_76[2],gpcOutL1_109[0],gpcOutL1_117[1],gpcOutL1_126[2]},gpcOutL2_51);
wire [2:0] gpcOutL2_52;

// (* RLOC = "X2Y52" *)
gpc006 gpcL2_52 ({gpcOutL1_57[0],gpcOutL1_63[1],gpcOutL1_69[2],gpcOutL1_101[0],gpcOutL1_109[1],gpcOutL1_117[2]},gpcOutL2_52);
wire [2:0] gpcOutL2_53;

// (* RLOC = "X2Y53" *)
gpc006 gpcL2_53 ({gpcOutL1_86[0],gpcOutL1_94[1],gpcOutL1_102[2],gpcOutL1_138[0],gpcOutL1_148[1],gpcOutL1_158[2]},gpcOutL2_53);
wire [2:0] gpcOutL2_54;

// (* RLOC = "X2Y54" *)
gpc006 gpcL2_54 ({gpcOutL1_65[0],gpcOutL1_71[1],gpcOutL1_78[2],gpcOutL1_111[0],gpcOutL1_119[1],gpcOutL1_128[2]},gpcOutL2_54);
wire [2:0] gpcOutL2_55;

// (* RLOC = "X2Y55" *)
gpc006 gpcL2_55 ({gpcOutL1_59[0],gpcOutL1_65[1],gpcOutL1_71[2],gpcOutL1_103[0],gpcOutL1_111[1],gpcOutL1_119[2]},gpcOutL2_55);
wire [2:0] gpcOutL2_56;

// (* RLOC = "X2Y56" *)
gpc006 gpcL2_56 ({gpcOutL1_92[0],gpcOutL1_100[1],gpcOutL1_108[2],gpcOutL1_146[0],gpcOutL1_156[1],gpcOutL1_166[2]},gpcOutL2_56);
wire [2:0] gpcOutL2_57;

// (* RLOC = "X2Y57" *)
gpc006 gpcL2_57 ({gpcOutL1_76[0],gpcOutL1_84[1],gpcOutL1_92[2],gpcOutL1_126[0],gpcOutL1_136[1],gpcOutL1_146[2]},gpcOutL2_57);
wire [2:0] gpcOutL2_58;

// (* RLOC = "X2Y58" *)
gpc006 gpcL2_58 ({gpcOutL1_94[0],gpcOutL1_102[1],gpcOutL1_110[2],gpcOutL1_148[0],gpcOutL1_158[1],gpcOutL1_168[2]},gpcOutL2_58);
wire [2:0] gpcOutL2_59;

// (* RLOC = "X2Y59" *)
gpc006 gpcL2_59 ({gpcOutL1_78[0],gpcOutL1_86[1],gpcOutL1_94[2],gpcOutL1_128[0],gpcOutL1_138[1],gpcOutL1_148[2]},gpcOutL2_59);
wire [2:0] gpcOutL2_60;

// (* RLOC = "X2Y60" *)
gpc006 gpcL2_60 ({gpcOutL1_81[2],gpcOutL1_89[1],gpcOutL1_97[0],gpcOutL1_131[2],gpcOutL1_141[1],gpcOutL1_151[0]},gpcOutL2_60);
wire [2:0] gpcOutL2_61;

// (* RLOC = "X2Y61" *)
gpc006 gpcL2_61 ({gpcOutL1_83[2],gpcOutL1_91[1],gpcOutL1_99[0],gpcOutL1_133[2],gpcOutL1_143[1],gpcOutL1_153[0]},gpcOutL2_61);
wire [2:0] gpcOutL2_62;

// (* RLOC = "X2Y62" *)
gpc006 gpcL2_62 ({gpcOutL1_116[0],gpcOutL1_125[1],gpcOutL1_135[2],gpcOutL1_176[0],gpcOutL1_187[1],gpcOutL1_199[2]},gpcOutL2_62);
wire [2:0] gpcOutL2_63;

// (* RLOC = "X2Y63" *)
gpc006 gpcL2_63 ({gpcOutL1_118[0],gpcOutL1_127[1],gpcOutL1_137[2],gpcOutL1_178[0],gpcOutL1_189[1],gpcOutL1_201[2]},gpcOutL2_63);
wire [2:0] gpcOutL2_64;

// (* RLOC = "X2Y64" *)
gpc006 gpcL2_64 ({gpcOutL1_89[2],gpcOutL1_97[1],gpcOutL1_105[0],gpcOutL1_141[2],gpcOutL1_151[1],gpcOutL1_161[0]},gpcOutL2_64);
wire [2:0] gpcOutL2_65;

// (* RLOC = "X2Y65" *)
gpc006 gpcL2_65 ({gpcOutL1_97[2],gpcOutL1_105[1],gpcOutL1_113[0],gpcOutL1_151[2],gpcOutL1_161[1],gpcOutL1_171[0]},gpcOutL2_65);
wire [2:0] gpcOutL2_66;

// (* RLOC = "X2Y66" *)
gpc006 gpcL2_66 ({gpcOutL1_105[2],gpcOutL1_113[1],gpcOutL1_122[0],gpcOutL1_161[2],gpcOutL1_171[1],gpcOutL1_182[0]},gpcOutL2_66);
wire [2:0] gpcOutL2_67;

// (* RLOC = "X2Y67" *)
gpc006 gpcL2_67 ({gpcOutL1_113[2],gpcOutL1_122[1],gpcOutL1_132[0],gpcOutL1_171[2],gpcOutL1_182[1],gpcOutL1_194[0]},gpcOutL2_67);
wire [2:0] gpcOutL2_68;

// (* RLOC = "X2Y68" *)
gpc006 gpcL2_68 ({gpcOutL1_122[2],gpcOutL1_132[1],gpcOutL1_142[0],gpcOutL1_182[2],gpcOutL1_194[1],gpcOutL1_206[0]},gpcOutL2_68);
wire [2:0] gpcOutL2_69;

// (* RLOC = "X2Y69" *)
gpc006 gpcL2_69 ({gpcOutL1_91[2],gpcOutL1_99[1],gpcOutL1_107[0],gpcOutL1_143[2],gpcOutL1_153[1],gpcOutL1_163[0]},gpcOutL2_69);
wire [2:0] gpcOutL2_70;

// (* RLOC = "X2Y70" *)
gpc006 gpcL2_70 ({gpcOutL1_99[2],gpcOutL1_107[1],gpcOutL1_115[0],gpcOutL1_153[2],gpcOutL1_163[1],gpcOutL1_173[0]},gpcOutL2_70);
wire [2:0] gpcOutL2_71;

// (* RLOC = "X2Y71" *)
gpc006 gpcL2_71 ({gpcOutL1_107[2],gpcOutL1_115[1],gpcOutL1_124[0],gpcOutL1_163[2],gpcOutL1_173[1],gpcOutL1_184[0]},gpcOutL2_71);
wire [2:0] gpcOutL2_72;

// (* RLOC = "X2Y72" *)
gpc006 gpcL2_72 ({gpcOutL1_115[2],gpcOutL1_124[1],gpcOutL1_134[0],gpcOutL1_173[2],gpcOutL1_184[1],gpcOutL1_196[0]},gpcOutL2_72);
wire [2:0] gpcOutL2_73;

// (* RLOC = "X2Y73" *)
gpc006 gpcL2_73 ({gpcOutL1_124[2],gpcOutL1_134[1],gpcOutL1_144[0],gpcOutL1_184[2],gpcOutL1_196[1],gpcOutL1_208[0]},gpcOutL2_73);
wire [2:0] gpcOutL2_74;

// (* RLOC = "X2Y74" *)
gpc006 gpcL2_74 ({gpcOutL1_135[0],gpcOutL1_145[1],gpcOutL1_155[2],gpcOutL1_199[0],gpcOutL1_211[1],gpcOutL1_223[2]},gpcOutL2_74);
wire [2:0] gpcOutL2_75;

// (* RLOC = "X2Y75" *)
gpc006 gpcL2_75 ({gpcOutL1_108[0],gpcOutL1_116[1],gpcOutL1_125[2],gpcOutL1_166[0],gpcOutL1_176[1],gpcOutL1_187[2]},gpcOutL2_75);
wire [2:0] gpcOutL2_76;

// (* RLOC = "X2Y76" *)
gpc006 gpcL2_76 ({gpcOutL1_100[0],gpcOutL1_108[1],gpcOutL1_116[2],gpcOutL1_156[0],gpcOutL1_166[1],gpcOutL1_176[2]},gpcOutL2_76);
wire [2:0] gpcOutL2_77;

// (* RLOC = "X2Y77" *)
gpc006 gpcL2_77 ({gpcOutL1_137[0],gpcOutL1_147[1],gpcOutL1_157[2],gpcOutL1_201[0],gpcOutL1_213[1],gpcOutL1_225[2]},gpcOutL2_77);
wire [2:0] gpcOutL2_78;

// (* RLOC = "X2Y78" *)
gpc006 gpcL2_78 ({gpcOutL1_110[0],gpcOutL1_118[1],gpcOutL1_127[2],gpcOutL1_168[0],gpcOutL1_178[1],gpcOutL1_189[2]},gpcOutL2_78);
wire [2:0] gpcOutL2_79;

// (* RLOC = "X2Y79" *)
gpc006 gpcL2_79 ({gpcOutL1_102[0],gpcOutL1_110[1],gpcOutL1_118[2],gpcOutL1_158[0],gpcOutL1_168[1],gpcOutL1_178[2]},gpcOutL2_79);
wire [2:0] gpcOutL2_80;

// (* RLOC = "X2Y80" *)
gpc006 gpcL2_80 ({gpcOutL1_139[0],gpcOutL1_149[1],gpcOutL1_159[2],gpcOutL1_203[0],gpcOutL1_215[1],gpcOutL1_227[2]},gpcOutL2_80);
wire [2:0] gpcOutL2_81;

// (* RLOC = "X2Y81" *)
gpc006 gpcL2_81 ({gpcOutL1_120[0],gpcOutL1_129[1],gpcOutL1_139[2],gpcOutL1_180[0],gpcOutL1_191[1],gpcOutL1_203[2]},gpcOutL2_81);
wire [2:0] gpcOutL2_82;

// (* RLOC = "X2Y82" *)
gpc006 gpcL2_82 ({gpcOutL1_120[1],gpcOutL1_129[2],gpcOutL1_130[0],gpcOutL1_180[1],gpcOutL1_191[2],gpcOutL1_192[0]},gpcOutL2_82);
wire [2:0] gpcOutL2_83;

// (* RLOC = "X2Y83" *)
gpc006 gpcL2_83 ({gpcOutL1_120[2],gpcOutL1_130[1],gpcOutL1_140[0],gpcOutL1_180[2],gpcOutL1_192[1],gpcOutL1_204[0]},gpcOutL2_83);
wire [2:0] gpcOutL2_84;

// (* RLOC = "X2Y84" *)
gpc006 gpcL2_84 ({gpcOutL1_130[2],gpcOutL1_140[1],gpcOutL1_150[0],gpcOutL1_192[2],gpcOutL1_204[1],gpcOutL1_216[0]},gpcOutL2_84);
wire [2:0] gpcOutL2_85;

// (* RLOC = "X2Y85" *)
gpc006 gpcL2_85 ({gpcOutL1_145[0],gpcOutL1_155[1],gpcOutL1_165[2],gpcOutL1_211[0],gpcOutL1_223[1],gpcOutL1_235[2]},gpcOutL2_85);
wire [2:0] gpcOutL2_86;

// (* RLOC = "X2Y86" *)
gpc006 gpcL2_86 ({gpcOutL1_125[0],gpcOutL1_135[1],gpcOutL1_145[2],gpcOutL1_187[0],gpcOutL1_199[1],gpcOutL1_211[2]},gpcOutL2_86);
wire [2:0] gpcOutL2_87;

// (* RLOC = "X2Y87" *)
gpc006 gpcL2_87 ({gpcOutL1_147[0],gpcOutL1_157[1],gpcOutL1_167[2],gpcOutL1_213[0],gpcOutL1_225[1],gpcOutL1_237[2]},gpcOutL2_87);
wire [2:0] gpcOutL2_88;

// (* RLOC = "X2Y88" *)
gpc006 gpcL2_88 ({gpcOutL1_127[0],gpcOutL1_137[1],gpcOutL1_147[2],gpcOutL1_189[0],gpcOutL1_201[1],gpcOutL1_213[2]},gpcOutL2_88);
wire [2:0] gpcOutL2_89;

// (* RLOC = "X2Y89" *)
gpc006 gpcL2_89 ({gpcOutL1_149[0],gpcOutL1_159[1],gpcOutL1_169[2],gpcOutL1_215[0],gpcOutL1_227[1],gpcOutL1_239[2]},gpcOutL2_89);
wire [2:0] gpcOutL2_90;

// (* RLOC = "X2Y90" *)
gpc006 gpcL2_90 ({gpcOutL1_129[0],gpcOutL1_139[1],gpcOutL1_149[2],gpcOutL1_191[0],gpcOutL1_203[1],gpcOutL1_215[2]},gpcOutL2_90);
wire [2:0] gpcOutL2_91;

// (* RLOC = "X2Y91" *)
gpc006 gpcL2_91 ({gpcOutL1_132[2],gpcOutL1_142[1],gpcOutL1_152[0],gpcOutL1_194[2],gpcOutL1_206[1],gpcOutL1_218[0]},gpcOutL2_91);
wire [2:0] gpcOutL2_92;

// (* RLOC = "X2Y92" *)
gpc006 gpcL2_92 ({gpcOutL1_134[2],gpcOutL1_144[1],gpcOutL1_154[0],gpcOutL1_196[2],gpcOutL1_208[1],gpcOutL1_220[0]},gpcOutL2_92);
wire [2:0] gpcOutL2_93;

// (* RLOC = "X2Y93" *)
gpc006 gpcL2_93 ({gpcOutL1_175[0],gpcOutL1_186[1],gpcOutL1_198[2],gpcOutL1_247[0],gpcOutL1_260[1],gpcOutL1_274[2]},gpcOutL2_93);
wire [2:0] gpcOutL2_94;

// (* RLOC = "X2Y94" *)
gpc006 gpcL2_94 ({gpcOutL1_177[0],gpcOutL1_188[1],gpcOutL1_200[2],gpcOutL1_249[0],gpcOutL1_262[1],gpcOutL1_276[2]},gpcOutL2_94);
wire [2:0] gpcOutL2_95;

// (* RLOC = "X2Y95" *)
gpc006 gpcL2_95 ({gpcOutL1_179[0],gpcOutL1_190[1],gpcOutL1_202[2],gpcOutL1_251[0],gpcOutL1_264[1],gpcOutL1_278[2]},gpcOutL2_95);
wire [2:0] gpcOutL2_96;

// (* RLOC = "X2Y96" *)
gpc006 gpcL2_96 ({gpcOutL1_140[2],gpcOutL1_150[1],gpcOutL1_160[0],gpcOutL1_204[2],gpcOutL1_216[1],gpcOutL1_228[0]},gpcOutL2_96);
wire [2:0] gpcOutL2_97;

// (* RLOC = "X2Y97" *)
gpc006 gpcL2_97 ({gpcOutL1_150[2],gpcOutL1_160[1],gpcOutL1_170[0],gpcOutL1_216[2],gpcOutL1_228[1],gpcOutL1_240[0]},gpcOutL2_97);
wire [2:0] gpcOutL2_98;

// (* RLOC = "X2Y98" *)
gpc006 gpcL2_98 ({gpcOutL1_160[2],gpcOutL1_170[1],gpcOutL1_181[0],gpcOutL1_228[2],gpcOutL1_240[1],gpcOutL1_253[0]},gpcOutL2_98);
wire [2:0] gpcOutL2_99;

// (* RLOC = "X2Y99" *)
gpc006 gpcL2_99 ({gpcOutL1_170[2],gpcOutL1_181[1],gpcOutL1_193[0],gpcOutL1_240[2],gpcOutL1_253[1],gpcOutL1_267[0]},gpcOutL2_99);
wire [2:0] gpcOutL2_100;

// (* RLOC = "X2Y100" *)
gpc006 gpcL2_100 ({gpcOutL1_181[2],gpcOutL1_193[1],gpcOutL1_205[0],gpcOutL1_253[2],gpcOutL1_267[1],gpcOutL1_281[0]},gpcOutL2_100);
wire [2:0] gpcOutL2_101;

// (* RLOC = "X2Y101" *)
gpc006 gpcL2_101 ({gpcOutL1_142[2],gpcOutL1_152[1],gpcOutL1_162[0],gpcOutL1_206[2],gpcOutL1_218[1],gpcOutL1_230[0]},gpcOutL2_101);
wire [2:0] gpcOutL2_102;

// (* RLOC = "X2Y102" *)
gpc006 gpcL2_102 ({gpcOutL1_152[2],gpcOutL1_162[1],gpcOutL1_172[0],gpcOutL1_218[2],gpcOutL1_230[1],gpcOutL1_242[0]},gpcOutL2_102);
wire [2:0] gpcOutL2_103;

// (* RLOC = "X2Y103" *)
gpc006 gpcL2_103 ({gpcOutL1_162[2],gpcOutL1_172[1],gpcOutL1_183[0],gpcOutL1_230[2],gpcOutL1_242[1],gpcOutL1_255[0]},gpcOutL2_103);
wire [2:0] gpcOutL2_104;

// (* RLOC = "X2Y104" *)
gpc006 gpcL2_104 ({gpcOutL1_172[2],gpcOutL1_183[1],gpcOutL1_195[0],gpcOutL1_242[2],gpcOutL1_255[1],gpcOutL1_269[0]},gpcOutL2_104);
wire [2:0] gpcOutL2_105;

// (* RLOC = "X2Y105" *)
gpc006 gpcL2_105 ({gpcOutL1_183[2],gpcOutL1_195[1],gpcOutL1_207[0],gpcOutL1_255[2],gpcOutL1_269[1],gpcOutL1_283[0]},gpcOutL2_105);
wire [2:0] gpcOutL2_106;

// (* RLOC = "X2Y106" *)
gpc006 gpcL2_106 ({gpcOutL1_144[2],gpcOutL1_154[1],gpcOutL1_164[0],gpcOutL1_208[2],gpcOutL1_220[1],gpcOutL1_232[0]},gpcOutL2_106);
wire [2:0] gpcOutL2_107;

// (* RLOC = "X2Y107" *)
gpc006 gpcL2_107 ({gpcOutL1_154[2],gpcOutL1_164[1],gpcOutL1_174[0],gpcOutL1_220[2],gpcOutL1_232[1],gpcOutL1_244[0]},gpcOutL2_107);
wire [2:0] gpcOutL2_108;

// (* RLOC = "X2Y108" *)
gpc006 gpcL2_108 ({gpcOutL1_164[2],gpcOutL1_174[1],gpcOutL1_185[0],gpcOutL1_232[2],gpcOutL1_244[1],gpcOutL1_257[0]},gpcOutL2_108);
wire [2:0] gpcOutL2_109;

// (* RLOC = "X2Y109" *)
gpc006 gpcL2_109 ({gpcOutL1_174[2],gpcOutL1_185[1],gpcOutL1_197[0],gpcOutL1_244[2],gpcOutL1_257[1],gpcOutL1_271[0]},gpcOutL2_109);
wire [2:0] gpcOutL2_110;

// (* RLOC = "X2Y110" *)
gpc006 gpcL2_110 ({gpcOutL1_185[2],gpcOutL1_197[1],gpcOutL1_209[0],gpcOutL1_257[2],gpcOutL1_271[1],gpcOutL1_285[0]},gpcOutL2_110);
wire [2:0] gpcOutL2_111;

// (* RLOC = "X2Y111" *)
gpc006 gpcL2_111 ({gpcOutL1_198[0],gpcOutL1_210[1],gpcOutL1_222[2],gpcOutL1_274[0],gpcOutL1_288[1],gpcOutL1_302[2]},gpcOutL2_111);
wire [2:0] gpcOutL2_112;

// (* RLOC = "X2Y112" *)
gpc006 gpcL2_112 ({gpcOutL1_165[0],gpcOutL1_175[1],gpcOutL1_186[2],gpcOutL1_235[0],gpcOutL1_247[1],gpcOutL1_260[2]},gpcOutL2_112);
wire [2:0] gpcOutL2_113;

// (* RLOC = "X2Y113" *)
gpc006 gpcL2_113 ({gpcOutL1_155[0],gpcOutL1_165[1],gpcOutL1_175[2],gpcOutL1_223[0],gpcOutL1_235[1],gpcOutL1_247[2]},gpcOutL2_113);
wire [2:0] gpcOutL2_114;

// (* RLOC = "X2Y114" *)
gpc006 gpcL2_114 ({gpcOutL1_200[0],gpcOutL1_212[1],gpcOutL1_224[2],gpcOutL1_276[0],gpcOutL1_290[1],gpcOutL1_304[2]},gpcOutL2_114);
wire [2:0] gpcOutL2_115;

// (* RLOC = "X2Y115" *)
gpc006 gpcL2_115 ({gpcOutL1_167[0],gpcOutL1_177[1],gpcOutL1_188[2],gpcOutL1_237[0],gpcOutL1_249[1],gpcOutL1_262[2]},gpcOutL2_115);
wire [2:0] gpcOutL2_116;

// (* RLOC = "X2Y116" *)
gpc006 gpcL2_116 ({gpcOutL1_157[0],gpcOutL1_167[1],gpcOutL1_177[2],gpcOutL1_225[0],gpcOutL1_237[1],gpcOutL1_249[2]},gpcOutL2_116);
wire [2:0] gpcOutL2_117;

// (* RLOC = "X2Y117" *)
gpc006 gpcL2_117 ({gpcOutL1_202[0],gpcOutL1_214[1],gpcOutL1_226[2],gpcOutL1_278[0],gpcOutL1_292[1],gpcOutL1_306[2]},gpcOutL2_117);
wire [2:0] gpcOutL2_118;

// (* RLOC = "X2Y118" *)
gpc006 gpcL2_118 ({gpcOutL1_169[0],gpcOutL1_179[1],gpcOutL1_190[2],gpcOutL1_239[0],gpcOutL1_251[1],gpcOutL1_264[2]},gpcOutL2_118);
wire [2:0] gpcOutL2_119;

// (* RLOC = "X2Y119" *)
gpc006 gpcL2_119 ({gpcOutL1_159[0],gpcOutL1_169[1],gpcOutL1_179[2],gpcOutL1_227[0],gpcOutL1_239[1],gpcOutL1_251[2]},gpcOutL2_119);
wire [2:0] gpcOutL2_120;

// (* RLOC = "X2Y120" *)
gpc006 gpcL2_120 ({gpcOutL1_210[0],gpcOutL1_222[1],gpcOutL1_234[2],gpcOutL1_288[0],gpcOutL1_302[1],gpcOutL1_316[2]},gpcOutL2_120);
wire [2:0] gpcOutL2_121;

// (* RLOC = "X2Y121" *)
gpc006 gpcL2_121 ({gpcOutL1_186[0],gpcOutL1_198[1],gpcOutL1_210[2],gpcOutL1_260[0],gpcOutL1_274[1],gpcOutL1_288[2]},gpcOutL2_121);
wire [2:0] gpcOutL2_122;

// (* RLOC = "X2Y122" *)
gpc006 gpcL2_122 ({gpcOutL1_212[0],gpcOutL1_224[1],gpcOutL1_236[2],gpcOutL1_290[0],gpcOutL1_304[1],gpcOutL1_318[2]},gpcOutL2_122);
wire [2:0] gpcOutL2_123;

// (* RLOC = "X2Y123" *)
gpc006 gpcL2_123 ({gpcOutL1_188[0],gpcOutL1_200[1],gpcOutL1_212[2],gpcOutL1_262[0],gpcOutL1_276[1],gpcOutL1_290[2]},gpcOutL2_123);
wire [2:0] gpcOutL2_124;

// (* RLOC = "X2Y124" *)
gpc006 gpcL2_124 ({gpcOutL1_214[0],gpcOutL1_226[1],gpcOutL1_238[2],gpcOutL1_292[0],gpcOutL1_306[1],gpcOutL1_320[2]},gpcOutL2_124);
wire [2:0] gpcOutL2_125;

// (* RLOC = "X2Y125" *)
gpc006 gpcL2_125 ({gpcOutL1_190[0],gpcOutL1_202[1],gpcOutL1_214[2],gpcOutL1_264[0],gpcOutL1_278[1],gpcOutL1_292[2]},gpcOutL2_125);
wire [2:0] gpcOutL2_126;

// (* RLOC = "X2Y126" *)
gpc006 gpcL2_126 ({gpcOutL1_193[2],gpcOutL1_205[1],gpcOutL1_217[0],gpcOutL1_267[2],gpcOutL1_281[1],gpcOutL1_295[0]},gpcOutL2_126);
wire [2:0] gpcOutL2_127;

// (* RLOC = "X2Y127" *)
gpc006 gpcL2_127 ({gpcOutL1_195[2],gpcOutL1_207[1],gpcOutL1_219[0],gpcOutL1_269[2],gpcOutL1_283[1],gpcOutL1_297[0]},gpcOutL2_127);
wire [2:0] gpcOutL2_128;

// (* RLOC = "X2Y128" *)
gpc006 gpcL2_128 ({gpcOutL1_197[2],gpcOutL1_209[1],gpcOutL1_221[0],gpcOutL1_271[2],gpcOutL1_285[1],gpcOutL1_299[0]},gpcOutL2_128);
wire [2:0] gpcOutL2_129;

// (* RLOC = "X2Y129" *)
gpc006 gpcL2_129 ({gpcOutL1_246[0],gpcOutL1_259[1],gpcOutL1_273[2],gpcOutL1_330[0],gpcOutL1_345[1],gpcOutL1_361[2]},gpcOutL2_129);
wire [2:0] gpcOutL2_130;

// (* RLOC = "X2Y130" *)
gpc006 gpcL2_130 ({gpcOutL1_248[0],gpcOutL1_261[1],gpcOutL1_275[2],gpcOutL1_332[0],gpcOutL1_347[1],gpcOutL1_363[2]},gpcOutL2_130);
wire [2:0] gpcOutL2_131;

// (* RLOC = "X2Y131" *)
gpc006 gpcL2_131 ({gpcOutL1_250[0],gpcOutL1_263[1],gpcOutL1_277[2],gpcOutL1_334[0],gpcOutL1_349[1],gpcOutL1_365[2]},gpcOutL2_131);
wire [2:0] gpcOutL2_132;

// (* RLOC = "X2Y132" *)
gpc006 gpcL2_132 ({gpcOutL1_205[2],gpcOutL1_217[1],gpcOutL1_229[0],gpcOutL1_281[2],gpcOutL1_295[1],gpcOutL1_309[0]},gpcOutL2_132);
wire [2:0] gpcOutL2_133;

// (* RLOC = "X2Y133" *)
gpc006 gpcL2_133 ({gpcOutL1_217[2],gpcOutL1_229[1],gpcOutL1_241[0],gpcOutL1_295[2],gpcOutL1_309[1],gpcOutL1_323[0]},gpcOutL2_133);
wire [2:0] gpcOutL2_134;

// (* RLOC = "X2Y134" *)
gpc006 gpcL2_134 ({gpcOutL1_229[2],gpcOutL1_241[1],gpcOutL1_254[0],gpcOutL1_309[2],gpcOutL1_323[1],gpcOutL1_338[0]},gpcOutL2_134);
wire [2:0] gpcOutL2_135;

// (* RLOC = "X2Y135" *)
gpc006 gpcL2_135 ({gpcOutL1_241[2],gpcOutL1_254[1],gpcOutL1_268[0],gpcOutL1_323[2],gpcOutL1_338[1],gpcOutL1_354[0]},gpcOutL2_135);
wire [2:0] gpcOutL2_136;

// (* RLOC = "X2Y136" *)
gpc006 gpcL2_136 ({gpcOutL1_254[2],gpcOutL1_268[1],gpcOutL1_282[0],gpcOutL1_338[2],gpcOutL1_354[1],gpcOutL1_370[0]},gpcOutL2_136);
wire [2:0] gpcOutL2_137;

// (* RLOC = "X2Y137" *)
gpc006 gpcL2_137 ({gpcOutL1_207[2],gpcOutL1_219[1],gpcOutL1_231[0],gpcOutL1_283[2],gpcOutL1_297[1],gpcOutL1_311[0]},gpcOutL2_137);
wire [2:0] gpcOutL2_138;

// (* RLOC = "X2Y138" *)
gpc006 gpcL2_138 ({gpcOutL1_219[2],gpcOutL1_231[1],gpcOutL1_243[0],gpcOutL1_297[2],gpcOutL1_311[1],gpcOutL1_325[0]},gpcOutL2_138);
wire [2:0] gpcOutL2_139;

// (* RLOC = "X2Y139" *)
gpc006 gpcL2_139 ({gpcOutL1_231[2],gpcOutL1_243[1],gpcOutL1_256[0],gpcOutL1_311[2],gpcOutL1_325[1],gpcOutL1_340[0]},gpcOutL2_139);
wire [2:0] gpcOutL2_140;

// (* RLOC = "X2Y140" *)
gpc006 gpcL2_140 ({gpcOutL1_243[2],gpcOutL1_256[1],gpcOutL1_270[0],gpcOutL1_325[2],gpcOutL1_340[1],gpcOutL1_356[0]},gpcOutL2_140);
wire [2:0] gpcOutL2_141;

// (* RLOC = "X2Y141" *)
gpc006 gpcL2_141 ({gpcOutL1_256[2],gpcOutL1_270[1],gpcOutL1_284[0],gpcOutL1_340[2],gpcOutL1_356[1],gpcOutL1_372[0]},gpcOutL2_141);
wire [2:0] gpcOutL2_142;

// (* RLOC = "X2Y142" *)
gpc006 gpcL2_142 ({gpcOutL1_209[2],gpcOutL1_221[1],gpcOutL1_233[0],gpcOutL1_285[2],gpcOutL1_299[1],gpcOutL1_313[0]},gpcOutL2_142);
wire [2:0] gpcOutL2_143;

// (* RLOC = "X2Y143" *)
gpc006 gpcL2_143 ({gpcOutL1_221[2],gpcOutL1_233[1],gpcOutL1_245[0],gpcOutL1_299[2],gpcOutL1_313[1],gpcOutL1_327[0]},gpcOutL2_143);
wire [2:0] gpcOutL2_144;

// (* RLOC = "X2Y144" *)
gpc006 gpcL2_144 ({gpcOutL1_233[2],gpcOutL1_245[1],gpcOutL1_258[0],gpcOutL1_313[2],gpcOutL1_327[1],gpcOutL1_342[0]},gpcOutL2_144);
wire [2:0] gpcOutL2_145;

// (* RLOC = "X2Y145" *)
gpc006 gpcL2_145 ({gpcOutL1_245[2],gpcOutL1_258[1],gpcOutL1_272[0],gpcOutL1_327[2],gpcOutL1_342[1],gpcOutL1_358[0]},gpcOutL2_145);
wire [2:0] gpcOutL2_146;

// (* RLOC = "X2Y146" *)
gpc006 gpcL2_146 ({gpcOutL1_258[2],gpcOutL1_272[1],gpcOutL1_286[0],gpcOutL1_342[2],gpcOutL1_358[1],gpcOutL1_374[0]},gpcOutL2_146);
wire [2:0] gpcOutL2_147;

// (* RLOC = "X2Y147" *)
gpc006 gpcL2_147 ({gpcOutL1_273[0],gpcOutL1_287[1],gpcOutL1_301[2],gpcOutL1_361[0],gpcOutL1_377[1],gpcOutL1_393[2]},gpcOutL2_147);
wire [2:0] gpcOutL2_148;

// (* RLOC = "X2Y148" *)
gpc006 gpcL2_148 ({gpcOutL1_234[0],gpcOutL1_246[1],gpcOutL1_259[2],gpcOutL1_316[0],gpcOutL1_330[1],gpcOutL1_345[2]},gpcOutL2_148);
wire [2:0] gpcOutL2_149;

// (* RLOC = "X2Y149" *)
gpc006 gpcL2_149 ({gpcOutL1_222[0],gpcOutL1_234[1],gpcOutL1_246[2],gpcOutL1_302[0],gpcOutL1_316[1],gpcOutL1_330[2]},gpcOutL2_149);
wire [2:0] gpcOutL2_150;

// (* RLOC = "X2Y150" *)
gpc006 gpcL2_150 ({gpcOutL1_275[0],gpcOutL1_289[1],gpcOutL1_303[2],gpcOutL1_363[0],gpcOutL1_379[1],gpcOutL1_395[2]},gpcOutL2_150);
wire [2:0] gpcOutL2_151;

// (* RLOC = "X2Y151" *)
gpc006 gpcL2_151 ({gpcOutL1_236[0],gpcOutL1_248[1],gpcOutL1_261[2],gpcOutL1_318[0],gpcOutL1_332[1],gpcOutL1_347[2]},gpcOutL2_151);
wire [2:0] gpcOutL2_152;

// (* RLOC = "X2Y152" *)
gpc006 gpcL2_152 ({gpcOutL1_224[0],gpcOutL1_236[1],gpcOutL1_248[2],gpcOutL1_304[0],gpcOutL1_318[1],gpcOutL1_332[2]},gpcOutL2_152);
wire [2:0] gpcOutL2_153;

// (* RLOC = "X2Y153" *)
gpc006 gpcL2_153 ({gpcOutL1_277[0],gpcOutL1_291[1],gpcOutL1_305[2],gpcOutL1_365[0],gpcOutL1_381[1],gpcOutL1_397[2]},gpcOutL2_153);
wire [2:0] gpcOutL2_154;

// (* RLOC = "X2Y154" *)
gpc006 gpcL2_154 ({gpcOutL1_238[0],gpcOutL1_250[1],gpcOutL1_263[2],gpcOutL1_320[0],gpcOutL1_334[1],gpcOutL1_349[2]},gpcOutL2_154);
wire [2:0] gpcOutL2_155;

// (* RLOC = "X2Y155" *)
gpc006 gpcL2_155 ({gpcOutL1_226[0],gpcOutL1_238[1],gpcOutL1_250[2],gpcOutL1_306[0],gpcOutL1_320[1],gpcOutL1_334[2]},gpcOutL2_155);
wire [2:0] gpcOutL2_156;

// (* RLOC = "X2Y156" *)
gpc006 gpcL2_156 ({gpcOutL1_279[0],gpcOutL1_293[1],gpcOutL1_307[2],gpcOutL1_367[0],gpcOutL1_383[1],gpcOutL1_399[2]},gpcOutL2_156);
wire [2:0] gpcOutL2_157;

// (* RLOC = "X2Y157" *)
gpc006 gpcL2_157 ({gpcOutL1_252[0],gpcOutL1_265[1],gpcOutL1_279[2],gpcOutL1_336[0],gpcOutL1_351[1],gpcOutL1_367[2]},gpcOutL2_157);
wire [2:0] gpcOutL2_158;

// (* RLOC = "X2Y158" *)
gpc006 gpcL2_158 ({gpcOutL1_252[1],gpcOutL1_265[2],gpcOutL1_266[0],gpcOutL1_336[1],gpcOutL1_351[2],gpcOutL1_352[0]},gpcOutL2_158);
wire [2:0] gpcOutL2_159;

// (* RLOC = "X2Y159" *)
gpc006 gpcL2_159 ({gpcOutL1_252[2],gpcOutL1_266[1],gpcOutL1_280[0],gpcOutL1_336[2],gpcOutL1_352[1],gpcOutL1_368[0]},gpcOutL2_159);
wire [2:0] gpcOutL2_160;

// (* RLOC = "X2Y160" *)
gpc006 gpcL2_160 ({gpcOutL1_266[2],gpcOutL1_280[1],gpcOutL1_294[0],gpcOutL1_352[2],gpcOutL1_368[1],gpcOutL1_384[0]},gpcOutL2_160);
wire [2:0] gpcOutL2_161;

// (* RLOC = "X2Y161" *)
gpc006 gpcL2_161 ({gpcOutL1_287[0],gpcOutL1_301[1],gpcOutL1_315[2],gpcOutL1_377[0],gpcOutL1_393[1],gpcOutL1_409[2]},gpcOutL2_161);
wire [2:0] gpcOutL2_162;

// (* RLOC = "X2Y162" *)
gpc006 gpcL2_162 ({gpcOutL1_259[0],gpcOutL1_273[1],gpcOutL1_287[2],gpcOutL1_345[0],gpcOutL1_361[1],gpcOutL1_377[2]},gpcOutL2_162);
wire [2:0] gpcOutL2_163;

// (* RLOC = "X2Y163" *)
gpc006 gpcL2_163 ({gpcOutL1_289[0],gpcOutL1_303[1],gpcOutL1_317[2],gpcOutL1_379[0],gpcOutL1_395[1],gpcOutL1_411[2]},gpcOutL2_163);
wire [2:0] gpcOutL2_164;

// (* RLOC = "X2Y164" *)
gpc006 gpcL2_164 ({gpcOutL1_261[0],gpcOutL1_275[1],gpcOutL1_289[2],gpcOutL1_347[0],gpcOutL1_363[1],gpcOutL1_379[2]},gpcOutL2_164);
wire [2:0] gpcOutL2_165;

// (* RLOC = "X2Y165" *)
gpc006 gpcL2_165 ({gpcOutL1_291[0],gpcOutL1_305[1],gpcOutL1_319[2],gpcOutL1_381[0],gpcOutL1_397[1],gpcOutL1_413[2]},gpcOutL2_165);
wire [2:0] gpcOutL2_166;

// (* RLOC = "X2Y166" *)
gpc006 gpcL2_166 ({gpcOutL1_263[0],gpcOutL1_277[1],gpcOutL1_291[2],gpcOutL1_349[0],gpcOutL1_365[1],gpcOutL1_381[2]},gpcOutL2_166);
wire [2:0] gpcOutL2_167;

// (* RLOC = "X2Y167" *)
gpc006 gpcL2_167 ({gpcOutL1_293[0],gpcOutL1_307[1],gpcOutL1_321[2],gpcOutL1_383[0],gpcOutL1_399[1],gpcOutL1_415[2]},gpcOutL2_167);
wire [2:0] gpcOutL2_168;

// (* RLOC = "X2Y168" *)
gpc006 gpcL2_168 ({gpcOutL1_265[0],gpcOutL1_279[1],gpcOutL1_293[2],gpcOutL1_351[0],gpcOutL1_367[1],gpcOutL1_383[2]},gpcOutL2_168);
wire [2:0] gpcOutL2_169;

// (* RLOC = "X2Y169" *)
gpc006 gpcL2_169 ({gpcOutL1_268[2],gpcOutL1_282[1],gpcOutL1_296[0],gpcOutL1_354[2],gpcOutL1_370[1],gpcOutL1_386[0]},gpcOutL2_169);
wire [2:0] gpcOutL2_170;

// (* RLOC = "X2Y170" *)
gpc006 gpcL2_170 ({gpcOutL1_270[2],gpcOutL1_284[1],gpcOutL1_298[0],gpcOutL1_356[2],gpcOutL1_372[1],gpcOutL1_388[0]},gpcOutL2_170);
wire [2:0] gpcOutL2_171;

// (* RLOC = "X2Y171" *)
gpc006 gpcL2_171 ({gpcOutL1_272[2],gpcOutL1_286[1],gpcOutL1_300[0],gpcOutL1_358[2],gpcOutL1_374[1],gpcOutL1_390[0]},gpcOutL2_171);
wire [2:0] gpcOutL2_172;

// (* RLOC = "X2Y172" *)
gpc006 gpcL2_172 ({gpcOutL1_329[0],gpcOutL1_344[1],gpcOutL1_360[2],gpcOutL1_425[0],gpcOutL1_442[1],gpcOutL1_460[2]},gpcOutL2_172);
wire [2:0] gpcOutL2_173;

// (* RLOC = "X2Y173" *)
gpc006 gpcL2_173 ({gpcOutL1_331[0],gpcOutL1_346[1],gpcOutL1_362[2],gpcOutL1_427[0],gpcOutL1_444[1],gpcOutL1_462[2]},gpcOutL2_173);
wire [2:0] gpcOutL2_174;

// (* RLOC = "X2Y174" *)
gpc006 gpcL2_174 ({gpcOutL1_333[0],gpcOutL1_348[1],gpcOutL1_364[2],gpcOutL1_429[0],gpcOutL1_446[1],gpcOutL1_464[2]},gpcOutL2_174);
wire [2:0] gpcOutL2_175;

// (* RLOC = "X2Y175" *)
gpc006 gpcL2_175 ({gpcOutL1_335[0],gpcOutL1_350[1],gpcOutL1_366[2],gpcOutL1_431[0],gpcOutL1_448[1],gpcOutL1_466[2]},gpcOutL2_175);
wire [2:0] gpcOutL2_176;

// (* RLOC = "X2Y176" *)
gpc006 gpcL2_176 ({gpcOutL1_280[2],gpcOutL1_294[1],gpcOutL1_308[0],gpcOutL1_368[2],gpcOutL1_384[1],gpcOutL1_400[0]},gpcOutL2_176);
wire [2:0] gpcOutL2_177;

// (* RLOC = "X2Y177" *)
gpc006 gpcL2_177 ({gpcOutL1_294[2],gpcOutL1_308[1],gpcOutL1_322[0],gpcOutL1_384[2],gpcOutL1_400[1],gpcOutL1_416[0]},gpcOutL2_177);
wire [2:0] gpcOutL2_178;

// (* RLOC = "X2Y178" *)
gpc006 gpcL2_178 ({gpcOutL1_308[2],gpcOutL1_322[1],gpcOutL1_337[0],gpcOutL1_400[2],gpcOutL1_416[1],gpcOutL1_433[0]},gpcOutL2_178);
wire [2:0] gpcOutL2_179;

// (* RLOC = "X2Y179" *)
gpc006 gpcL2_179 ({gpcOutL1_322[2],gpcOutL1_337[1],gpcOutL1_353[0],gpcOutL1_416[2],gpcOutL1_433[1],gpcOutL1_451[0]},gpcOutL2_179);
wire [2:0] gpcOutL2_180;

// (* RLOC = "X2Y180" *)
gpc006 gpcL2_180 ({gpcOutL1_337[2],gpcOutL1_353[1],gpcOutL1_369[0],gpcOutL1_433[2],gpcOutL1_451[1],gpcOutL1_469[0]},gpcOutL2_180);
wire [2:0] gpcOutL2_181;

// (* RLOC = "X2Y181" *)
gpc006 gpcL2_181 ({gpcOutL1_282[2],gpcOutL1_296[1],gpcOutL1_310[0],gpcOutL1_370[2],gpcOutL1_386[1],gpcOutL1_402[0]},gpcOutL2_181);
wire [2:0] gpcOutL2_182;

// (* RLOC = "X2Y182" *)
gpc006 gpcL2_182 ({gpcOutL1_296[2],gpcOutL1_310[1],gpcOutL1_324[0],gpcOutL1_386[2],gpcOutL1_402[1],gpcOutL1_418[0]},gpcOutL2_182);
wire [2:0] gpcOutL2_183;

// (* RLOC = "X2Y183" *)
gpc006 gpcL2_183 ({gpcOutL1_310[2],gpcOutL1_324[1],gpcOutL1_339[0],gpcOutL1_402[2],gpcOutL1_418[1],gpcOutL1_435[0]},gpcOutL2_183);
wire [2:0] gpcOutL2_184;

// (* RLOC = "X2Y184" *)
gpc006 gpcL2_184 ({gpcOutL1_324[2],gpcOutL1_339[1],gpcOutL1_355[0],gpcOutL1_418[2],gpcOutL1_435[1],gpcOutL1_453[0]},gpcOutL2_184);
wire [2:0] gpcOutL2_185;

// (* RLOC = "X2Y185" *)
gpc006 gpcL2_185 ({gpcOutL1_339[2],gpcOutL1_355[1],gpcOutL1_371[0],gpcOutL1_435[2],gpcOutL1_453[1],gpcOutL1_471[0]},gpcOutL2_185);
wire [2:0] gpcOutL2_186;

// (* RLOC = "X2Y186" *)
gpc006 gpcL2_186 ({gpcOutL1_284[2],gpcOutL1_298[1],gpcOutL1_312[0],gpcOutL1_372[2],gpcOutL1_388[1],gpcOutL1_404[0]},gpcOutL2_186);
wire [2:0] gpcOutL2_187;

// (* RLOC = "X2Y187" *)
gpc006 gpcL2_187 ({gpcOutL1_298[2],gpcOutL1_312[1],gpcOutL1_326[0],gpcOutL1_388[2],gpcOutL1_404[1],gpcOutL1_420[0]},gpcOutL2_187);
wire [2:0] gpcOutL2_188;

// (* RLOC = "X2Y188" *)
gpc006 gpcL2_188 ({gpcOutL1_312[2],gpcOutL1_326[1],gpcOutL1_341[0],gpcOutL1_404[2],gpcOutL1_420[1],gpcOutL1_437[0]},gpcOutL2_188);
wire [2:0] gpcOutL2_189;

// (* RLOC = "X2Y189" *)
gpc006 gpcL2_189 ({gpcOutL1_326[2],gpcOutL1_341[1],gpcOutL1_357[0],gpcOutL1_420[2],gpcOutL1_437[1],gpcOutL1_455[0]},gpcOutL2_189);
wire [2:0] gpcOutL2_190;

// (* RLOC = "X2Y190" *)
gpc006 gpcL2_190 ({gpcOutL1_341[2],gpcOutL1_357[1],gpcOutL1_373[0],gpcOutL1_437[2],gpcOutL1_455[1],gpcOutL1_473[0]},gpcOutL2_190);
wire [2:0] gpcOutL2_191;

// (* RLOC = "X2Y191" *)
gpc006 gpcL2_191 ({gpcOutL1_286[2],gpcOutL1_300[1],gpcOutL1_314[0],gpcOutL1_374[2],gpcOutL1_390[1],gpcOutL1_406[0]},gpcOutL2_191);
wire [2:0] gpcOutL2_192;

// (* RLOC = "X2Y192" *)
gpc006 gpcL2_192 ({gpcOutL1_300[2],gpcOutL1_314[1],gpcOutL1_328[0],gpcOutL1_390[2],gpcOutL1_406[1],gpcOutL1_422[0]},gpcOutL2_192);
wire [2:0] gpcOutL2_193;

// (* RLOC = "X2Y193" *)
gpc006 gpcL2_193 ({gpcOutL1_314[2],gpcOutL1_328[1],gpcOutL1_343[0],gpcOutL1_406[2],gpcOutL1_422[1],gpcOutL1_439[0]},gpcOutL2_193);
wire [2:0] gpcOutL2_194;

// (* RLOC = "X2Y194" *)
gpc006 gpcL2_194 ({gpcOutL1_328[2],gpcOutL1_343[1],gpcOutL1_359[0],gpcOutL1_422[2],gpcOutL1_439[1],gpcOutL1_457[0]},gpcOutL2_194);
wire [2:0] gpcOutL2_195;

// (* RLOC = "X2Y195" *)
gpc006 gpcL2_195 ({gpcOutL1_343[2],gpcOutL1_359[1],gpcOutL1_375[0],gpcOutL1_439[2],gpcOutL1_457[1],gpcOutL1_475[0]},gpcOutL2_195);
wire [2:0] gpcOutL2_196;

// (* RLOC = "X2Y196" *)
gpc006 gpcL2_196 ({gpcOutL1_360[0],gpcOutL1_376[1],gpcOutL1_392[2],gpcOutL1_460[0],gpcOutL1_478[1],gpcOutL1_496[2]},gpcOutL2_196);
wire [2:0] gpcOutL2_197;

// (* RLOC = "X2Y197" *)
gpc006 gpcL2_197 ({gpcOutL1_315[0],gpcOutL1_329[1],gpcOutL1_344[2],gpcOutL1_409[0],gpcOutL1_425[1],gpcOutL1_442[2]},gpcOutL2_197);
wire [2:0] gpcOutL2_198;

// (* RLOC = "X2Y198" *)
gpc006 gpcL2_198 ({gpcOutL1_301[0],gpcOutL1_315[1],gpcOutL1_329[2],gpcOutL1_393[0],gpcOutL1_409[1],gpcOutL1_425[2]},gpcOutL2_198);
wire [2:0] gpcOutL2_199;

// (* RLOC = "X2Y199" *)
gpc006 gpcL2_199 ({gpcOutL1_362[0],gpcOutL1_378[1],gpcOutL1_394[2],gpcOutL1_462[0],gpcOutL1_480[1],gpcOutL1_498[2]},gpcOutL2_199);
wire [2:0] gpcOutL2_200;

// (* RLOC = "X2Y200" *)
gpc006 gpcL2_200 ({gpcOutL1_317[0],gpcOutL1_331[1],gpcOutL1_346[2],gpcOutL1_411[0],gpcOutL1_427[1],gpcOutL1_444[2]},gpcOutL2_200);
wire [2:0] gpcOutL2_201;

// (* RLOC = "X2Y201" *)
gpc006 gpcL2_201 ({gpcOutL1_303[0],gpcOutL1_317[1],gpcOutL1_331[2],gpcOutL1_395[0],gpcOutL1_411[1],gpcOutL1_427[2]},gpcOutL2_201);
wire [2:0] gpcOutL2_202;

// (* RLOC = "X2Y202" *)
gpc006 gpcL2_202 ({gpcOutL1_364[0],gpcOutL1_380[1],gpcOutL1_396[2],gpcOutL1_464[0],gpcOutL1_482[1],gpcOutL1_500[2]},gpcOutL2_202);
wire [2:0] gpcOutL2_203;

// (* RLOC = "X2Y203" *)
gpc006 gpcL2_203 ({gpcOutL1_319[0],gpcOutL1_333[1],gpcOutL1_348[2],gpcOutL1_413[0],gpcOutL1_429[1],gpcOutL1_446[2]},gpcOutL2_203);
wire [2:0] gpcOutL2_204;

// (* RLOC = "X2Y204" *)
gpc006 gpcL2_204 ({gpcOutL1_305[0],gpcOutL1_319[1],gpcOutL1_333[2],gpcOutL1_397[0],gpcOutL1_413[1],gpcOutL1_429[2]},gpcOutL2_204);
wire [2:0] gpcOutL2_205;

// (* RLOC = "X2Y205" *)
gpc006 gpcL2_205 ({gpcOutL1_366[0],gpcOutL1_382[1],gpcOutL1_398[2],gpcOutL1_466[0],gpcOutL1_484[1],gpcOutL1_502[2]},gpcOutL2_205);
wire [2:0] gpcOutL2_206;

// (* RLOC = "X2Y206" *)
gpc006 gpcL2_206 ({gpcOutL1_321[0],gpcOutL1_335[1],gpcOutL1_350[2],gpcOutL1_415[0],gpcOutL1_431[1],gpcOutL1_448[2]},gpcOutL2_206);
wire [2:0] gpcOutL2_207;

// (* RLOC = "X2Y207" *)
gpc006 gpcL2_207 ({gpcOutL1_307[0],gpcOutL1_321[1],gpcOutL1_335[2],gpcOutL1_399[0],gpcOutL1_415[1],gpcOutL1_431[2]},gpcOutL2_207);
wire [2:0] gpcOutL2_208;

// (* RLOC = "X2Y208" *)
gpc006 gpcL2_208 ({gpcOutL1_376[0],gpcOutL1_392[1],gpcOutL1_408[2],gpcOutL1_478[0],gpcOutL1_496[1],gpcOutL1_514[2]},gpcOutL2_208);
wire [2:0] gpcOutL2_209;

// (* RLOC = "X2Y209" *)
gpc006 gpcL2_209 ({gpcOutL1_344[0],gpcOutL1_360[1],gpcOutL1_376[2],gpcOutL1_442[0],gpcOutL1_460[1],gpcOutL1_478[2]},gpcOutL2_209);
wire [2:0] gpcOutL2_210;

// (* RLOC = "X2Y210" *)
gpc006 gpcL2_210 ({gpcOutL1_378[0],gpcOutL1_394[1],gpcOutL1_410[2],gpcOutL1_480[0],gpcOutL1_498[1],gpcOutL1_516[2]},gpcOutL2_210);
wire [2:0] gpcOutL2_211;

// (* RLOC = "X2Y211" *)
gpc006 gpcL2_211 ({gpcOutL1_346[0],gpcOutL1_362[1],gpcOutL1_378[2],gpcOutL1_444[0],gpcOutL1_462[1],gpcOutL1_480[2]},gpcOutL2_211);
wire [2:0] gpcOutL2_212;

// (* RLOC = "X2Y212" *)
gpc006 gpcL2_212 ({gpcOutL1_380[0],gpcOutL1_396[1],gpcOutL1_412[2],gpcOutL1_482[0],gpcOutL1_500[1],gpcOutL1_518[2]},gpcOutL2_212);
wire [2:0] gpcOutL2_213;

// (* RLOC = "X2Y213" *)
gpc006 gpcL2_213 ({gpcOutL1_348[0],gpcOutL1_364[1],gpcOutL1_380[2],gpcOutL1_446[0],gpcOutL1_464[1],gpcOutL1_482[2]},gpcOutL2_213);
wire [2:0] gpcOutL2_214;

// (* RLOC = "X2Y214" *)
gpc006 gpcL2_214 ({gpcOutL1_382[0],gpcOutL1_398[1],gpcOutL1_414[2],gpcOutL1_484[0],gpcOutL1_502[1],gpcOutL1_520[2]},gpcOutL2_214);
wire [2:0] gpcOutL2_215;

// (* RLOC = "X2Y215" *)
gpc006 gpcL2_215 ({gpcOutL1_350[0],gpcOutL1_366[1],gpcOutL1_382[2],gpcOutL1_448[0],gpcOutL1_466[1],gpcOutL1_484[2]},gpcOutL2_215);
wire [2:0] gpcOutL2_216;

// (* RLOC = "X2Y216" *)
gpc006 gpcL2_216 ({gpcOutL1_353[2],gpcOutL1_369[1],gpcOutL1_385[0],gpcOutL1_451[2],gpcOutL1_469[1],gpcOutL1_487[0]},gpcOutL2_216);
wire [2:0] gpcOutL2_217;

// (* RLOC = "X2Y217" *)
gpc006 gpcL2_217 ({gpcOutL1_355[2],gpcOutL1_371[1],gpcOutL1_387[0],gpcOutL1_453[2],gpcOutL1_471[1],gpcOutL1_489[0]},gpcOutL2_217);
wire [2:0] gpcOutL2_218;

// (* RLOC = "X2Y218" *)
gpc006 gpcL2_218 ({gpcOutL1_357[2],gpcOutL1_373[1],gpcOutL1_389[0],gpcOutL1_455[2],gpcOutL1_473[1],gpcOutL1_491[0]},gpcOutL2_218);
wire [2:0] gpcOutL2_219;

// (* RLOC = "X2Y219" *)
gpc006 gpcL2_219 ({gpcOutL1_359[2],gpcOutL1_375[1],gpcOutL1_391[0],gpcOutL1_457[2],gpcOutL1_475[1],gpcOutL1_493[0]},gpcOutL2_219);
wire [2:0] gpcOutL2_220;

// (* RLOC = "X2Y220" *)
gpc006 gpcL2_220 ({gpcOutL1_424[0],gpcOutL1_441[1],gpcOutL1_459[2],gpcOutL1_532[0],gpcOutL1_551[1],gpcOutL1_571[2]},gpcOutL2_220);
wire [2:0] gpcOutL2_221;

// (* RLOC = "X2Y221" *)
gpc006 gpcL2_221 ({gpcOutL1_426[0],gpcOutL1_443[1],gpcOutL1_461[2],gpcOutL1_534[0],gpcOutL1_553[1],gpcOutL1_573[2]},gpcOutL2_221);
wire [2:0] gpcOutL2_222;

// (* RLOC = "X2Y222" *)
gpc006 gpcL2_222 ({gpcOutL1_428[0],gpcOutL1_445[1],gpcOutL1_463[2],gpcOutL1_536[0],gpcOutL1_555[1],gpcOutL1_575[2]},gpcOutL2_222);
wire [2:0] gpcOutL2_223;

// (* RLOC = "X2Y223" *)
gpc006 gpcL2_223 ({gpcOutL1_430[0],gpcOutL1_447[1],gpcOutL1_465[2],gpcOutL1_538[0],gpcOutL1_557[1],gpcOutL1_577[2]},gpcOutL2_223);
wire [2:0] gpcOutL2_224;

// (* RLOC = "X2Y224" *)
gpc006 gpcL2_224 ({gpcOutL1_369[2],gpcOutL1_385[1],gpcOutL1_401[0],gpcOutL1_469[2],gpcOutL1_487[1],gpcOutL1_505[0]},gpcOutL2_224);
wire [2:0] gpcOutL2_225;

// (* RLOC = "X2Y225" *)
gpc006 gpcL2_225 ({gpcOutL1_385[2],gpcOutL1_401[1],gpcOutL1_417[0],gpcOutL1_487[2],gpcOutL1_505[1],gpcOutL1_523[0]},gpcOutL2_225);
wire [2:0] gpcOutL2_226;

// (* RLOC = "X2Y226" *)
gpc006 gpcL2_226 ({gpcOutL1_401[2],gpcOutL1_417[1],gpcOutL1_434[0],gpcOutL1_505[2],gpcOutL1_523[1],gpcOutL1_542[0]},gpcOutL2_226);
wire [2:0] gpcOutL2_227;

// (* RLOC = "X2Y227" *)
gpc006 gpcL2_227 ({gpcOutL1_417[2],gpcOutL1_434[1],gpcOutL1_452[0],gpcOutL1_523[2],gpcOutL1_542[1],gpcOutL1_562[0]},gpcOutL2_227);
wire [2:0] gpcOutL2_228;

// (* RLOC = "X2Y228" *)
gpc006 gpcL2_228 ({gpcOutL1_434[2],gpcOutL1_452[1],gpcOutL1_470[0],gpcOutL1_542[2],gpcOutL1_562[1],gpcOutL1_582[0]},gpcOutL2_228);
wire [2:0] gpcOutL2_229;

// (* RLOC = "X2Y229" *)
gpc006 gpcL2_229 ({gpcOutL1_371[2],gpcOutL1_387[1],gpcOutL1_403[0],gpcOutL1_471[2],gpcOutL1_489[1],gpcOutL1_507[0]},gpcOutL2_229);
wire [2:0] gpcOutL2_230;

// (* RLOC = "X2Y230" *)
gpc006 gpcL2_230 ({gpcOutL1_387[2],gpcOutL1_403[1],gpcOutL1_419[0],gpcOutL1_489[2],gpcOutL1_507[1],gpcOutL1_525[0]},gpcOutL2_230);
wire [2:0] gpcOutL2_231;

// (* RLOC = "X2Y231" *)
gpc006 gpcL2_231 ({gpcOutL1_403[2],gpcOutL1_419[1],gpcOutL1_436[0],gpcOutL1_507[2],gpcOutL1_525[1],gpcOutL1_544[0]},gpcOutL2_231);
wire [2:0] gpcOutL2_232;

// (* RLOC = "X2Y232" *)
gpc006 gpcL2_232 ({gpcOutL1_419[2],gpcOutL1_436[1],gpcOutL1_454[0],gpcOutL1_525[2],gpcOutL1_544[1],gpcOutL1_564[0]},gpcOutL2_232);
wire [2:0] gpcOutL2_233;

// (* RLOC = "X2Y233" *)
gpc006 gpcL2_233 ({gpcOutL1_436[2],gpcOutL1_454[1],gpcOutL1_472[0],gpcOutL1_544[2],gpcOutL1_564[1],gpcOutL1_584[0]},gpcOutL2_233);
wire [2:0] gpcOutL2_234;

// (* RLOC = "X2Y234" *)
gpc006 gpcL2_234 ({gpcOutL1_373[2],gpcOutL1_389[1],gpcOutL1_405[0],gpcOutL1_473[2],gpcOutL1_491[1],gpcOutL1_509[0]},gpcOutL2_234);
wire [2:0] gpcOutL2_235;

// (* RLOC = "X2Y235" *)
gpc006 gpcL2_235 ({gpcOutL1_389[2],gpcOutL1_405[1],gpcOutL1_421[0],gpcOutL1_491[2],gpcOutL1_509[1],gpcOutL1_527[0]},gpcOutL2_235);
wire [2:0] gpcOutL2_236;

// (* RLOC = "X2Y236" *)
gpc006 gpcL2_236 ({gpcOutL1_405[2],gpcOutL1_421[1],gpcOutL1_438[0],gpcOutL1_509[2],gpcOutL1_527[1],gpcOutL1_546[0]},gpcOutL2_236);
wire [2:0] gpcOutL2_237;

// (* RLOC = "X2Y237" *)
gpc006 gpcL2_237 ({gpcOutL1_421[2],gpcOutL1_438[1],gpcOutL1_456[0],gpcOutL1_527[2],gpcOutL1_546[1],gpcOutL1_566[0]},gpcOutL2_237);
wire [2:0] gpcOutL2_238;

// (* RLOC = "X2Y238" *)
gpc006 gpcL2_238 ({gpcOutL1_438[2],gpcOutL1_456[1],gpcOutL1_474[0],gpcOutL1_546[2],gpcOutL1_566[1],gpcOutL1_586[0]},gpcOutL2_238);
wire [2:0] gpcOutL2_239;

// (* RLOC = "X2Y239" *)
gpc006 gpcL2_239 ({gpcOutL1_375[2],gpcOutL1_391[1],gpcOutL1_407[0],gpcOutL1_475[2],gpcOutL1_493[1],gpcOutL1_511[0]},gpcOutL2_239);
wire [2:0] gpcOutL2_240;

// (* RLOC = "X2Y240" *)
gpc006 gpcL2_240 ({gpcOutL1_391[2],gpcOutL1_407[1],gpcOutL1_423[0],gpcOutL1_493[2],gpcOutL1_511[1],gpcOutL1_529[0]},gpcOutL2_240);
wire [2:0] gpcOutL2_241;

// (* RLOC = "X2Y241" *)
gpc006 gpcL2_241 ({gpcOutL1_407[2],gpcOutL1_423[1],gpcOutL1_440[0],gpcOutL1_511[2],gpcOutL1_529[1],gpcOutL1_548[0]},gpcOutL2_241);
wire [2:0] gpcOutL2_242;

// (* RLOC = "X2Y242" *)
gpc006 gpcL2_242 ({gpcOutL1_423[2],gpcOutL1_440[1],gpcOutL1_458[0],gpcOutL1_529[2],gpcOutL1_548[1],gpcOutL1_568[0]},gpcOutL2_242);
wire [2:0] gpcOutL2_243;

// (* RLOC = "X2Y243" *)
gpc006 gpcL2_243 ({gpcOutL1_440[2],gpcOutL1_458[1],gpcOutL1_476[0],gpcOutL1_548[2],gpcOutL1_568[1],gpcOutL1_588[0]},gpcOutL2_243);
wire [2:0] gpcOutL2_244;

// (* RLOC = "X2Y244" *)
gpc006 gpcL2_244 ({gpcOutL1_459[0],gpcOutL1_477[1],gpcOutL1_495[2],gpcOutL1_571[0],gpcOutL1_591[1],gpcOutL1_611[2]},gpcOutL2_244);
wire [2:0] gpcOutL2_245;

// (* RLOC = "X2Y245" *)
gpc006 gpcL2_245 ({gpcOutL1_408[0],gpcOutL1_424[1],gpcOutL1_441[2],gpcOutL1_514[0],gpcOutL1_532[1],gpcOutL1_551[2]},gpcOutL2_245);
wire [2:0] gpcOutL2_246;

// (* RLOC = "X2Y246" *)
gpc006 gpcL2_246 ({gpcOutL1_392[0],gpcOutL1_408[1],gpcOutL1_424[2],gpcOutL1_496[0],gpcOutL1_514[1],gpcOutL1_532[2]},gpcOutL2_246);
wire [2:0] gpcOutL2_247;

// (* RLOC = "X2Y247" *)
gpc006 gpcL2_247 ({gpcOutL1_461[0],gpcOutL1_479[1],gpcOutL1_497[2],gpcOutL1_573[0],gpcOutL1_593[1],gpcOutL1_613[2]},gpcOutL2_247);
wire [2:0] gpcOutL2_248;

// (* RLOC = "X2Y248" *)
gpc006 gpcL2_248 ({gpcOutL1_410[0],gpcOutL1_426[1],gpcOutL1_443[2],gpcOutL1_516[0],gpcOutL1_534[1],gpcOutL1_553[2]},gpcOutL2_248);
wire [2:0] gpcOutL2_249;

// (* RLOC = "X2Y249" *)
gpc006 gpcL2_249 ({gpcOutL1_394[0],gpcOutL1_410[1],gpcOutL1_426[2],gpcOutL1_498[0],gpcOutL1_516[1],gpcOutL1_534[2]},gpcOutL2_249);
wire [2:0] gpcOutL2_250;

// (* RLOC = "X2Y250" *)
gpc006 gpcL2_250 ({gpcOutL1_463[0],gpcOutL1_481[1],gpcOutL1_499[2],gpcOutL1_575[0],gpcOutL1_595[1],gpcOutL1_615[2]},gpcOutL2_250);
wire [2:0] gpcOutL2_251;

// (* RLOC = "X2Y251" *)
gpc006 gpcL2_251 ({gpcOutL1_412[0],gpcOutL1_428[1],gpcOutL1_445[2],gpcOutL1_518[0],gpcOutL1_536[1],gpcOutL1_555[2]},gpcOutL2_251);
wire [2:0] gpcOutL2_252;

// (* RLOC = "X2Y252" *)
gpc006 gpcL2_252 ({gpcOutL1_396[0],gpcOutL1_412[1],gpcOutL1_428[2],gpcOutL1_500[0],gpcOutL1_518[1],gpcOutL1_536[2]},gpcOutL2_252);
wire [2:0] gpcOutL2_253;

// (* RLOC = "X2Y253" *)
gpc006 gpcL2_253 ({gpcOutL1_465[0],gpcOutL1_483[1],gpcOutL1_501[2],gpcOutL1_577[0],gpcOutL1_597[1],gpcOutL1_617[2]},gpcOutL2_253);
wire [2:0] gpcOutL2_254;

// (* RLOC = "X2Y254" *)
gpc006 gpcL2_254 ({gpcOutL1_414[0],gpcOutL1_430[1],gpcOutL1_447[2],gpcOutL1_520[0],gpcOutL1_538[1],gpcOutL1_557[2]},gpcOutL2_254);
wire [2:0] gpcOutL2_255;

// (* RLOC = "X2Y255" *)
gpc006 gpcL2_255 ({gpcOutL1_398[0],gpcOutL1_414[1],gpcOutL1_430[2],gpcOutL1_502[0],gpcOutL1_520[1],gpcOutL1_538[2]},gpcOutL2_255);
wire [2:0] gpcOutL2_256;

// (* RLOC = "X2Y256" *)
gpc006 gpcL2_256 ({gpcOutL1_467[0],gpcOutL1_485[1],gpcOutL1_503[2],gpcOutL1_579[0],gpcOutL1_599[1],gpcOutL1_619[2]},gpcOutL2_256);
wire [2:0] gpcOutL2_257;

// (* RLOC = "X2Y257" *)
gpc006 gpcL2_257 ({gpcOutL1_432[0],gpcOutL1_449[1],gpcOutL1_467[2],gpcOutL1_540[0],gpcOutL1_559[1],gpcOutL1_579[2]},gpcOutL2_257);
wire [2:0] gpcOutL2_258;

// (* RLOC = "X2Y258" *)
gpc006 gpcL2_258 ({gpcOutL1_432[1],gpcOutL1_449[2],gpcOutL1_450[0],gpcOutL1_540[1],gpcOutL1_559[2],gpcOutL1_560[0]},gpcOutL2_258);
wire [2:0] gpcOutL2_259;

// (* RLOC = "X2Y259" *)
gpc006 gpcL2_259 ({gpcOutL1_432[2],gpcOutL1_450[1],gpcOutL1_468[0],gpcOutL1_540[2],gpcOutL1_560[1],gpcOutL1_580[0]},gpcOutL2_259);
wire [2:0] gpcOutL2_260;

// (* RLOC = "X2Y260" *)
gpc006 gpcL2_260 ({gpcOutL1_450[2],gpcOutL1_468[1],gpcOutL1_486[0],gpcOutL1_560[2],gpcOutL1_580[1],gpcOutL1_600[0]},gpcOutL2_260);
wire [2:0] gpcOutL2_261;

// (* RLOC = "X2Y261" *)
gpc006 gpcL2_261 ({gpcOutL1_477[0],gpcOutL1_495[1],gpcOutL1_513[2],gpcOutL1_591[0],gpcOutL1_611[1],gpcOutL1_631[2]},gpcOutL2_261);
wire [2:0] gpcOutL2_262;

// (* RLOC = "X2Y262" *)
gpc006 gpcL2_262 ({gpcOutL1_441[0],gpcOutL1_459[1],gpcOutL1_477[2],gpcOutL1_551[0],gpcOutL1_571[1],gpcOutL1_591[2]},gpcOutL2_262);
wire [2:0] gpcOutL2_263;

// (* RLOC = "X2Y263" *)
gpc006 gpcL2_263 ({gpcOutL1_479[0],gpcOutL1_497[1],gpcOutL1_515[2],gpcOutL1_593[0],gpcOutL1_613[1],gpcOutL1_633[2]},gpcOutL2_263);
wire [2:0] gpcOutL2_264;

// (* RLOC = "X2Y264" *)
gpc006 gpcL2_264 ({gpcOutL1_443[0],gpcOutL1_461[1],gpcOutL1_479[2],gpcOutL1_553[0],gpcOutL1_573[1],gpcOutL1_593[2]},gpcOutL2_264);
wire [2:0] gpcOutL2_265;

// (* RLOC = "X2Y265" *)
gpc006 gpcL2_265 ({gpcOutL1_481[0],gpcOutL1_499[1],gpcOutL1_517[2],gpcOutL1_595[0],gpcOutL1_615[1],gpcOutL1_635[2]},gpcOutL2_265);
wire [2:0] gpcOutL2_266;

// (* RLOC = "X2Y266" *)
gpc006 gpcL2_266 ({gpcOutL1_445[0],gpcOutL1_463[1],gpcOutL1_481[2],gpcOutL1_555[0],gpcOutL1_575[1],gpcOutL1_595[2]},gpcOutL2_266);
wire [2:0] gpcOutL2_267;

// (* RLOC = "X2Y267" *)
gpc006 gpcL2_267 ({gpcOutL1_483[0],gpcOutL1_501[1],gpcOutL1_519[2],gpcOutL1_597[0],gpcOutL1_617[1],gpcOutL1_637[2]},gpcOutL2_267);
wire [2:0] gpcOutL2_268;

// (* RLOC = "X2Y268" *)
gpc006 gpcL2_268 ({gpcOutL1_447[0],gpcOutL1_465[1],gpcOutL1_483[2],gpcOutL1_557[0],gpcOutL1_577[1],gpcOutL1_597[2]},gpcOutL2_268);
wire [2:0] gpcOutL2_269;

// (* RLOC = "X2Y269" *)
gpc006 gpcL2_269 ({gpcOutL1_485[0],gpcOutL1_503[1],gpcOutL1_521[2],gpcOutL1_599[0],gpcOutL1_619[1],gpcOutL1_639[2]},gpcOutL2_269);
wire [2:0] gpcOutL2_270;

// (* RLOC = "X2Y270" *)
gpc006 gpcL2_270 ({gpcOutL1_449[0],gpcOutL1_467[1],gpcOutL1_485[2],gpcOutL1_559[0],gpcOutL1_579[1],gpcOutL1_599[2]},gpcOutL2_270);
wire [2:0] gpcOutL2_271;

// (* RLOC = "X2Y271" *)
gpc006 gpcL2_271 ({gpcOutL1_452[2],gpcOutL1_470[1],gpcOutL1_488[0],gpcOutL1_562[2],gpcOutL1_582[1],gpcOutL1_602[0]},gpcOutL2_271);
wire [2:0] gpcOutL2_272;

// (* RLOC = "X2Y272" *)
gpc006 gpcL2_272 ({gpcOutL1_454[2],gpcOutL1_472[1],gpcOutL1_490[0],gpcOutL1_564[2],gpcOutL1_584[1],gpcOutL1_604[0]},gpcOutL2_272);
wire [2:0] gpcOutL2_273;

// (* RLOC = "X2Y273" *)
gpc006 gpcL2_273 ({gpcOutL1_456[2],gpcOutL1_474[1],gpcOutL1_492[0],gpcOutL1_566[2],gpcOutL1_586[1],gpcOutL1_606[0]},gpcOutL2_273);
wire [2:0] gpcOutL2_274;

// (* RLOC = "X2Y274" *)
gpc006 gpcL2_274 ({gpcOutL1_458[2],gpcOutL1_476[1],gpcOutL1_494[0],gpcOutL1_568[2],gpcOutL1_588[1],gpcOutL1_608[0]},gpcOutL2_274);
wire [2:0] gpcOutL2_275;

// (* RLOC = "X2Y275" *)
gpc006 gpcL2_275 ({gpcOutL1_531[0],gpcOutL1_550[1],gpcOutL1_570[2],gpcOutL1_651[1],pp8[1],pp9[0]},gpcOutL2_275);
wire [2:0] gpcOutL2_276;

// (* RLOC = "X2Y276" *)
gpc006 gpcL2_276 ({gpcOutL1_533[0],gpcOutL1_552[1],gpcOutL1_572[2],gpcOutL1_653[1],pp20[1],pp21[0]},gpcOutL2_276);
wire [2:0] gpcOutL2_277;

// (* RLOC = "X2Y277" *)
gpc006 gpcL2_277 ({gpcOutL1_535[0],gpcOutL1_554[1],gpcOutL1_574[2],gpcOutL1_655[1],pp32[1],pp33[0]},gpcOutL2_277);
wire [2:0] gpcOutL2_278;

// (* RLOC = "X2Y278" *)
gpc006 gpcL2_278 ({gpcOutL1_537[0],gpcOutL1_556[1],gpcOutL1_576[2],gpcOutL1_657[1],pp44[1],pp45[0]},gpcOutL2_278);
wire [2:0] gpcOutL2_279;

// (* RLOC = "X2Y279" *)
gpc006 gpcL2_279 ({gpcOutL1_539[0],gpcOutL1_558[1],gpcOutL1_578[2],gpcOutL1_659[1],pp56[1],pp57[0]},gpcOutL2_279);
wire [2:0] gpcOutL2_280;

// (* RLOC = "X2Y280" *)
gpc006 gpcL2_280 ({gpcOutL1_468[2],gpcOutL1_486[1],gpcOutL1_504[0],gpcOutL1_580[2],gpcOutL1_600[1],gpcOutL1_620[0]},gpcOutL2_280);
wire [2:0] gpcOutL2_281;

// (* RLOC = "X2Y281" *)
gpc006 gpcL2_281 ({gpcOutL1_486[2],gpcOutL1_504[1],gpcOutL1_522[0],gpcOutL1_600[2],gpcOutL1_620[1],gpcOutL1_640[0]},gpcOutL2_281);
wire [2:0] gpcOutL2_282;

// (* RLOC = "X2Y282" *)
gpc006 gpcL2_282 ({gpcOutL1_504[2],gpcOutL1_522[1],gpcOutL1_541[0],gpcOutL1_620[2],gpcOutL1_640[1],gpcOutL1_662[0]},gpcOutL2_282);
wire [2:0] gpcOutL2_283;

// (* RLOC = "X2Y283" *)
gpc006 gpcL2_283 ({gpcOutL1_522[2],gpcOutL1_541[1],gpcOutL1_561[0],gpcOutL1_640[2],gpcOutL1_662[1],pp63[7]},gpcOutL2_283);
wire [2:0] gpcOutL2_284;

// (* RLOC = "X2Y284" *)
gpc006 gpcL2_284 ({gpcOutL1_541[2],gpcOutL1_561[1],gpcOutL1_581[0],gpcOutL1_662[2],pp62[9],pp63[8]},gpcOutL2_284);
wire [2:0] gpcOutL2_285;

// (* RLOC = "X2Y285" *)
gpc006 gpcL2_285 ({gpcOutL1_470[2],gpcOutL1_488[1],gpcOutL1_506[0],gpcOutL1_582[2],gpcOutL1_602[1],gpcOutL1_622[0]},gpcOutL2_285);
wire [2:0] gpcOutL2_286;

// (* RLOC = "X2Y286" *)
gpc006 gpcL2_286 ({gpcOutL1_488[2],gpcOutL1_506[1],gpcOutL1_524[0],gpcOutL1_602[2],gpcOutL1_622[1],gpcOutL1_642[0]},gpcOutL2_286);
wire [2:0] gpcOutL2_287;

// (* RLOC = "X2Y287" *)
gpc006 gpcL2_287 ({gpcOutL1_506[2],gpcOutL1_524[1],gpcOutL1_543[0],gpcOutL1_622[2],gpcOutL1_642[1],gpcOutL1_664[0]},gpcOutL2_287);
wire [2:0] gpcOutL2_288;

// (* RLOC = "X2Y288" *)
gpc006 gpcL2_288 ({gpcOutL1_524[2],gpcOutL1_543[1],gpcOutL1_563[0],gpcOutL1_642[2],gpcOutL1_664[1],pp63[19]},gpcOutL2_288);
wire [2:0] gpcOutL2_289;

// (* RLOC = "X2Y289" *)
gpc006 gpcL2_289 ({gpcOutL1_543[2],gpcOutL1_563[1],gpcOutL1_583[0],gpcOutL1_664[2],pp62[21],pp63[20]},gpcOutL2_289);
wire [2:0] gpcOutL2_290;

// (* RLOC = "X2Y290" *)
gpc006 gpcL2_290 ({gpcOutL1_472[2],gpcOutL1_490[1],gpcOutL1_508[0],gpcOutL1_584[2],gpcOutL1_604[1],gpcOutL1_624[0]},gpcOutL2_290);
wire [2:0] gpcOutL2_291;

// (* RLOC = "X2Y291" *)
gpc006 gpcL2_291 ({gpcOutL1_490[2],gpcOutL1_508[1],gpcOutL1_526[0],gpcOutL1_604[2],gpcOutL1_624[1],gpcOutL1_644[0]},gpcOutL2_291);
wire [2:0] gpcOutL2_292;

// (* RLOC = "X2Y292" *)
gpc006 gpcL2_292 ({gpcOutL1_508[2],gpcOutL1_526[1],gpcOutL1_545[0],gpcOutL1_624[2],gpcOutL1_644[1],gpcOutL1_666[0]},gpcOutL2_292);
wire [2:0] gpcOutL2_293;

// (* RLOC = "X2Y293" *)
gpc006 gpcL2_293 ({gpcOutL1_526[2],gpcOutL1_545[1],gpcOutL1_565[0],gpcOutL1_644[2],gpcOutL1_666[1],pp63[31]},gpcOutL2_293);
wire [2:0] gpcOutL2_294;

// (* RLOC = "X2Y294" *)
gpc006 gpcL2_294 ({gpcOutL1_545[2],gpcOutL1_565[1],gpcOutL1_585[0],gpcOutL1_666[2],pp62[33],pp63[32]},gpcOutL2_294);
wire [2:0] gpcOutL2_295;

// (* RLOC = "X2Y295" *)
gpc006 gpcL2_295 ({gpcOutL1_474[2],gpcOutL1_492[1],gpcOutL1_510[0],gpcOutL1_586[2],gpcOutL1_606[1],gpcOutL1_626[0]},gpcOutL2_295);
wire [2:0] gpcOutL2_296;

// (* RLOC = "X2Y296" *)
gpc006 gpcL2_296 ({gpcOutL1_492[2],gpcOutL1_510[1],gpcOutL1_528[0],gpcOutL1_606[2],gpcOutL1_626[1],gpcOutL1_646[0]},gpcOutL2_296);
wire [2:0] gpcOutL2_297;

// (* RLOC = "X2Y297" *)
gpc006 gpcL2_297 ({gpcOutL1_510[2],gpcOutL1_528[1],gpcOutL1_547[0],gpcOutL1_626[2],gpcOutL1_646[1],gpcOutL1_668[0]},gpcOutL2_297);
wire [2:0] gpcOutL2_298;

// (* RLOC = "X2Y298" *)
gpc006 gpcL2_298 ({gpcOutL1_528[2],gpcOutL1_547[1],gpcOutL1_567[0],gpcOutL1_646[2],gpcOutL1_668[1],pp63[43]},gpcOutL2_298);
wire [2:0] gpcOutL2_299;

// (* RLOC = "X2Y299" *)
gpc006 gpcL2_299 ({gpcOutL1_547[2],gpcOutL1_567[1],gpcOutL1_587[0],gpcOutL1_668[2],pp62[45],pp63[44]},gpcOutL2_299);
wire [2:0] gpcOutL2_300;

// (* RLOC = "X2Y300" *)
gpc006 gpcL2_300 ({gpcOutL1_476[2],gpcOutL1_494[1],gpcOutL1_512[0],gpcOutL1_588[2],gpcOutL1_608[1],gpcOutL1_628[0]},gpcOutL2_300);
wire [2:0] gpcOutL2_301;

// (* RLOC = "X2Y301" *)
gpc006 gpcL2_301 ({gpcOutL1_494[2],gpcOutL1_512[1],gpcOutL1_530[0],gpcOutL1_608[2],gpcOutL1_628[1],gpcOutL1_648[0]},gpcOutL2_301);
wire [2:0] gpcOutL2_302;

// (* RLOC = "X2Y302" *)
gpc006 gpcL2_302 ({gpcOutL1_512[2],gpcOutL1_530[1],gpcOutL1_549[0],gpcOutL1_628[2],gpcOutL1_648[1],gpcOutL1_670[0]},gpcOutL2_302);
wire [2:0] gpcOutL2_303;

// (* RLOC = "X2Y303" *)
gpc006 gpcL2_303 ({gpcOutL1_530[2],gpcOutL1_549[1],gpcOutL1_569[0],gpcOutL1_648[2],gpcOutL1_670[1],pp63[55]},gpcOutL2_303);
wire [2:0] gpcOutL2_304;

// (* RLOC = "X2Y304" *)
gpc006 gpcL2_304 ({gpcOutL1_549[2],gpcOutL1_569[1],gpcOutL1_589[0],gpcOutL1_670[2],pp62[57],pp63[56]},gpcOutL2_304);
wire [2:0] gpcOutL2_305;

// (* RLOC = "X2Y305" *)
gpc015 gpcL2_305 ({gpcOutL1_550[0],gpcOutL1_570[0],gpcOutL1_590[1],gpcOutL1_610[2],pp6[1],pp7[0]},gpcOutL2_305);
wire [2:0] gpcOutL2_306;

// (* RLOC = "X2Y306" *)
gpc015 gpcL2_306 ({gpcOutL1_495[0],gpcOutL1_513[0],gpcOutL1_531[1],gpcOutL1_550[2],gpcOutL1_631[0],gpcOutL1_651[2]},gpcOutL2_306);
wire [2:0] gpcOutL2_307;

// (* RLOC = "X2Y307" *)
gpc015 gpcL2_307 ({gpcOutL1_552[0],gpcOutL1_572[0],gpcOutL1_592[1],gpcOutL1_612[2],pp18[1],pp19[0]},gpcOutL2_307);
wire [2:0] gpcOutL2_308;

// (* RLOC = "X2Y308" *)
gpc015 gpcL2_308 ({gpcOutL1_497[0],gpcOutL1_515[0],gpcOutL1_533[1],gpcOutL1_552[2],gpcOutL1_633[0],gpcOutL1_653[2]},gpcOutL2_308);
wire [2:0] gpcOutL2_309;

// (* RLOC = "X2Y309" *)
gpc015 gpcL2_309 ({gpcOutL1_554[0],gpcOutL1_574[0],gpcOutL1_594[1],gpcOutL1_614[2],pp30[1],pp31[0]},gpcOutL2_309);
wire [2:0] gpcOutL2_310;

// (* RLOC = "X2Y310" *)
gpc015 gpcL2_310 ({gpcOutL1_499[0],gpcOutL1_517[0],gpcOutL1_535[1],gpcOutL1_554[2],gpcOutL1_635[0],gpcOutL1_655[2]},gpcOutL2_310);
wire [2:0] gpcOutL2_311;

// (* RLOC = "X2Y311" *)
gpc015 gpcL2_311 ({gpcOutL1_556[0],gpcOutL1_576[0],gpcOutL1_596[1],gpcOutL1_616[2],pp42[1],pp43[0]},gpcOutL2_311);
wire [2:0] gpcOutL2_312;

// (* RLOC = "X2Y312" *)
gpc015 gpcL2_312 ({gpcOutL1_501[0],gpcOutL1_519[0],gpcOutL1_537[1],gpcOutL1_556[2],gpcOutL1_637[0],gpcOutL1_657[2]},gpcOutL2_312);
wire [2:0] gpcOutL2_313;

// (* RLOC = "X2Y313" *)
gpc015 gpcL2_313 ({gpcOutL1_558[0],gpcOutL1_578[0],gpcOutL1_598[1],gpcOutL1_618[2],pp54[1],pp55[0]},gpcOutL2_313);
wire [2:0] gpcOutL2_314;

// (* RLOC = "X2Y314" *)
gpc015 gpcL2_314 ({gpcOutL1_503[0],gpcOutL1_521[0],gpcOutL1_539[1],gpcOutL1_558[2],gpcOutL1_639[0],gpcOutL1_659[2]},gpcOutL2_314);
wire [3:0] gpcOutL2_315;

// (* RLOC = "X2Y315" *)
gpc042 gpcL2_315 ({gpcOutL1_590[0],gpcOutL1_610[1],gpcOutL1_630[2],pp6[0],gpcOutL1_610[0],gpcOutL1_630[1]},gpcOutL2_315);
wire [2:0] gpcOutL2_316;

// (* RLOC = "X2Y316" *)
gpc014 gpcL2_316 ({pp12[0],gpcOutL1_513[1],gpcOutL1_531[2],gpcOutL1_611[0],gpcOutL1_631[1]},gpcOutL2_316);
wire [3:0] gpcOutL2_317;

// (* RLOC = "X2Y317" *)
gpc042 gpcL2_317 ({gpcOutL1_592[0],gpcOutL1_612[1],gpcOutL1_632[2],pp18[0],gpcOutL1_612[0],gpcOutL1_632[1]},gpcOutL2_317);
wire [2:0] gpcOutL2_318;

// (* RLOC = "X2Y318" *)
gpc014 gpcL2_318 ({pp24[0],gpcOutL1_515[1],gpcOutL1_533[2],gpcOutL1_613[0],gpcOutL1_633[1]},gpcOutL2_318);
wire [3:0] gpcOutL2_319;

// (* RLOC = "X2Y319" *)
gpc042 gpcL2_319 ({gpcOutL1_594[0],gpcOutL1_614[1],gpcOutL1_634[2],pp30[0],gpcOutL1_614[0],gpcOutL1_634[1]},gpcOutL2_319);
wire [2:0] gpcOutL2_320;

// (* RLOC = "X2Y320" *)
gpc014 gpcL2_320 ({pp36[0],gpcOutL1_517[1],gpcOutL1_535[2],gpcOutL1_615[0],gpcOutL1_635[1]},gpcOutL2_320);
wire [3:0] gpcOutL2_321;

// (* RLOC = "X2Y321" *)
gpc042 gpcL2_321 ({gpcOutL1_596[0],gpcOutL1_616[1],gpcOutL1_636[2],pp42[0],gpcOutL1_616[0],gpcOutL1_636[1]},gpcOutL2_321);
wire [2:0] gpcOutL2_322;

// (* RLOC = "X2Y322" *)
gpc014 gpcL2_322 ({pp48[0],gpcOutL1_519[1],gpcOutL1_537[2],gpcOutL1_617[0],gpcOutL1_637[1]},gpcOutL2_322);
wire [3:0] gpcOutL2_323;

// (* RLOC = "X2Y323" *)
gpc042 gpcL2_323 ({gpcOutL1_598[0],gpcOutL1_618[1],gpcOutL1_638[2],pp54[0],gpcOutL1_618[0],gpcOutL1_638[1]},gpcOutL2_323);
wire [2:0] gpcOutL2_324;

// (* RLOC = "X2Y324" *)
gpc014 gpcL2_324 ({pp60[0],gpcOutL1_521[1],gpcOutL1_539[2],gpcOutL1_619[0],gpcOutL1_639[1]},gpcOutL2_324);
wire [2:0] gpcOutL2_325;

// (* RLOC = "X2Y325" *)
gpc014 gpcL2_325 ({gpcOutL1_581[2],gpcOutL1_561[2],gpcOutL1_581[1],gpcOutL1_601[0],pp63[9]},gpcOutL2_325);
wire [2:0] gpcOutL2_326;

// (* RLOC = "X2Y326" *)
gpc014 gpcL2_326 ({gpcOutL1_583[2],gpcOutL1_563[2],gpcOutL1_583[1],gpcOutL1_603[0],pp63[21]},gpcOutL2_326);
wire [2:0] gpcOutL2_327;

// (* RLOC = "X2Y327" *)
gpc014 gpcL2_327 ({gpcOutL1_585[2],gpcOutL1_565[2],gpcOutL1_585[1],gpcOutL1_605[0],pp63[33]},gpcOutL2_327);
wire [2:0] gpcOutL2_328;

// (* RLOC = "X2Y328" *)
gpc014 gpcL2_328 ({gpcOutL1_587[2],gpcOutL1_567[2],gpcOutL1_587[1],gpcOutL1_607[0],pp63[45]},gpcOutL2_328);
wire [2:0] gpcOutL2_329;

// (* RLOC = "X2Y329" *)
gpc014 gpcL2_329 ({gpcOutL1_589[2],gpcOutL1_569[2],gpcOutL1_589[1],gpcOutL1_609[0],pp63[57]},gpcOutL2_329);
wire [2:0] gpcOutL2_330;

// (* RLOC = "X2Y330" *)
gpc023 gpcL2_330 ({gpcOutL1_630[0],gpcOutL1_650[2],gpcOutL1_650[1],pp2[1],pp3[0]},gpcOutL2_330);
wire [1:0] gpcOutL2_331;

// (* RLOC = "X2Y331" *)
gpc003 gpcL2_331 ({gpcOutL1_570[1],gpcOutL1_590[2],gpcOutL1_651[0]},gpcOutL2_331);
wire [2:0] gpcOutL2_332;

// (* RLOC = "X2Y332" *)
gpc023 gpcL2_332 ({gpcOutL1_632[0],gpcOutL1_652[2],gpcOutL1_652[1],pp14[1],pp15[0]},gpcOutL2_332);
wire [1:0] gpcOutL2_333;

// (* RLOC = "X2Y333" *)
gpc003 gpcL2_333 ({gpcOutL1_572[1],gpcOutL1_592[2],gpcOutL1_653[0]},gpcOutL2_333);
wire [2:0] gpcOutL2_334;

// (* RLOC = "X2Y334" *)
gpc023 gpcL2_334 ({gpcOutL1_634[0],gpcOutL1_654[2],gpcOutL1_654[1],pp26[1],pp27[0]},gpcOutL2_334);
wire [1:0] gpcOutL2_335;

// (* RLOC = "X2Y335" *)
gpc003 gpcL2_335 ({gpcOutL1_574[1],gpcOutL1_594[2],gpcOutL1_655[0]},gpcOutL2_335);
wire [2:0] gpcOutL2_336;

// (* RLOC = "X2Y336" *)
gpc023 gpcL2_336 ({gpcOutL1_636[0],gpcOutL1_656[2],gpcOutL1_656[1],pp38[1],pp39[0]},gpcOutL2_336);
wire [1:0] gpcOutL2_337;

// (* RLOC = "X2Y337" *)
gpc003 gpcL2_337 ({gpcOutL1_576[1],gpcOutL1_596[2],gpcOutL1_657[0]},gpcOutL2_337);
wire [2:0] gpcOutL2_338;

// (* RLOC = "X2Y338" *)
gpc023 gpcL2_338 ({gpcOutL1_638[0],gpcOutL1_658[2],gpcOutL1_658[1],pp50[1],pp51[0]},gpcOutL2_338);
wire [1:0] gpcOutL2_339;

// (* RLOC = "X2Y339" *)
gpc003 gpcL2_339 ({gpcOutL1_578[1],gpcOutL1_598[2],gpcOutL1_659[0]},gpcOutL2_339);
wire [2:0] gpcOutL2_340;

// (* RLOC = "X2Y340" *)
gpc023 gpcL2_340 ({gpcOutL1_621[2],gpcOutL1_641[1],gpcOutL1_601[2],gpcOutL1_621[1],gpcOutL1_641[0]},gpcOutL2_340);
wire [2:0] gpcOutL2_341;

// (* RLOC = "X2Y341" *)
gpc023 gpcL2_341 ({gpcOutL1_663[2],pp62[15],gpcOutL1_641[2],gpcOutL1_663[1],pp63[13]},gpcOutL2_341);
wire [2:0] gpcOutL2_342;

// (* RLOC = "X2Y342" *)
gpc023 gpcL2_342 ({gpcOutL1_623[2],gpcOutL1_643[1],gpcOutL1_603[2],gpcOutL1_623[1],gpcOutL1_643[0]},gpcOutL2_342);
wire [2:0] gpcOutL2_343;

// (* RLOC = "X2Y343" *)
gpc023 gpcL2_343 ({gpcOutL1_665[2],pp62[27],gpcOutL1_643[2],gpcOutL1_665[1],pp63[25]},gpcOutL2_343);
wire [2:0] gpcOutL2_344;

// (* RLOC = "X2Y344" *)
gpc023 gpcL2_344 ({gpcOutL1_625[2],gpcOutL1_645[1],gpcOutL1_605[2],gpcOutL1_625[1],gpcOutL1_645[0]},gpcOutL2_344);
wire [2:0] gpcOutL2_345;

// (* RLOC = "X2Y345" *)
gpc023 gpcL2_345 ({gpcOutL1_667[2],pp62[39],gpcOutL1_645[2],gpcOutL1_667[1],pp63[37]},gpcOutL2_345);
wire [2:0] gpcOutL2_346;

// (* RLOC = "X2Y346" *)
gpc023 gpcL2_346 ({gpcOutL1_627[2],gpcOutL1_647[1],gpcOutL1_607[2],gpcOutL1_627[1],gpcOutL1_647[0]},gpcOutL2_346);
wire [2:0] gpcOutL2_347;

// (* RLOC = "X2Y347" *)
gpc023 gpcL2_347 ({gpcOutL1_669[2],pp62[51],gpcOutL1_647[2],gpcOutL1_669[1],pp63[49]},gpcOutL2_347);
wire [2:0] gpcOutL2_348;

// (* RLOC = "X2Y348" *)
gpc023 gpcL2_348 ({gpcOutL1_629[2],gpcOutL1_649[1],gpcOutL1_609[2],gpcOutL1_629[1],gpcOutL1_649[0]},gpcOutL2_348);
wire [2:0] gpcOutL2_349;

// (* RLOC = "X2Y349" *)
gpc023 gpcL2_349 ({gpcOutL1_671[2],pp62[63],gpcOutL1_649[2],gpcOutL1_671[1],pp63[61]},gpcOutL2_349);
wire [3:0] gpcOutL2_350;

// (* RLOC = "X2Y350" *)
gpc212 gpcL2_350 ({gpcOutL1_660[0],gpcOutL1_661[1],gpcOutL1_661[0],pp60[1],pp61[0]},gpcOutL2_350);
wire [3:0] gpcOutL2_351;

// (* RLOC = "X2Y351" *)
gpc222 gpcL2_351 ({gpcOutL1_672[2],pp63[3],gpcOutL1_660[2],gpcOutL1_672[1],gpcOutL1_660[1],gpcOutL1_672[0]},gpcOutL2_351);
wire [2:0] gpcOutL3_0;

// (* RLOC = "X3Y0" *)
gpc006 gpcL3_0 ({gpcOutL2_1[1],gpcOutL2_2[0],gpcOutL2_6[2],gpcOutL2_29[1],gpcOutL2_30[0],gpcOutL2_36[2]},gpcOutL3_0);
wire [2:0] gpcOutL3_1;

// (* RLOC = "X3Y1" *)
gpc006 gpcL3_1 ({gpcOutL2_0[0],gpcOutL2_5[1],gpcOutL2_15[2],gpcOutL2_28[0],gpcOutL2_35[1],gpcOutL2_55[2]},gpcOutL3_1);
wire [2:0] gpcOutL3_2;

// (* RLOC = "X3Y2" *)
gpc006 gpcL3_2 ({gpcOutL2_0[1],gpcOutL2_5[2],gpcOutL2_6[0],gpcOutL2_28[1],gpcOutL2_35[2],gpcOutL2_36[0]},gpcOutL3_2);
wire [2:0] gpcOutL3_3;

// (* RLOC = "X3Y3" *)
gpc006 gpcL3_3 ({gpcOutL2_0[2],gpcOutL2_1[0],gpcOutL2_6[1],gpcOutL2_28[2],gpcOutL2_29[0],gpcOutL2_36[1]},gpcOutL3_3);
wire [2:0] gpcOutL3_4;

// (* RLOC = "X3Y4" *)
gpc006 gpcL3_4 ({gpcOutL2_1[2],gpcOutL2_2[1],gpcOutL2_3[0],gpcOutL2_29[2],gpcOutL2_30[1],gpcOutL2_31[0]},gpcOutL3_4);
wire [2:0] gpcOutL3_5;

// (* RLOC = "X3Y5" *)
gpc006 gpcL3_5 ({gpcOutL2_2[2],gpcOutL2_3[1],gpcOutL2_4[0],gpcOutL2_30[2],gpcOutL2_31[1],gpcOutL2_32[0]},gpcOutL3_5);
wire [2:0] gpcOutL3_6;

// (* RLOC = "X3Y6" *)
gpc006 gpcL3_6 ({gpcOutL2_3[2],gpcOutL2_4[1],gpcOutL2_8[0],gpcOutL2_31[2],gpcOutL2_32[1],gpcOutL2_40[0]},gpcOutL3_6);
wire [2:0] gpcOutL3_7;

// (* RLOC = "X3Y7" *)
gpc006 gpcL3_7 ({gpcOutL2_12[2],gpcOutL2_18[1],gpcOutL2_20[0],gpcOutL2_44[2],gpcOutL2_60[1],gpcOutL2_64[0]},gpcOutL3_7);
wire [2:0] gpcOutL3_8;

// (* RLOC = "X3Y8" *)
gpc006 gpcL3_8 ({gpcOutL2_13[1],gpcOutL2_16[2],gpcOutL2_17[0],gpcOutL2_53[1],gpcOutL2_58[2],gpcOutL2_59[0]},gpcOutL3_8);
wire [2:0] gpcOutL3_9;

// (* RLOC = "X3Y9" *)
gpc006 gpcL3_9 ({gpcOutL2_7[0],gpcOutL2_13[2],gpcOutL2_17[1],gpcOutL2_39[0],gpcOutL2_53[2],gpcOutL2_59[1]},gpcOutL3_9);
wire [2:0] gpcOutL3_10;

// (* RLOC = "X3Y10" *)
gpc006 gpcL3_10 ({gpcOutL2_7[2],gpcOutL2_14[1],gpcOutL2_15[0],gpcOutL2_39[2],gpcOutL2_54[1],gpcOutL2_55[0]},gpcOutL3_10);
wire [2:0] gpcOutL3_11;

// (* RLOC = "X3Y11" *)
gpc006 gpcL3_11 ({gpcOutL2_5[0],gpcOutL2_14[2],gpcOutL2_15[1],gpcOutL2_35[0],gpcOutL2_54[2],gpcOutL2_55[1]},gpcOutL3_11);
wire [2:0] gpcOutL3_12;

// (* RLOC = "X3Y12" *)
gpc006 gpcL3_12 ({gpcOutL2_4[2],gpcOutL2_8[1],gpcOutL2_9[0],gpcOutL2_32[2],gpcOutL2_40[1],gpcOutL2_41[0]},gpcOutL3_12);
wire [2:0] gpcOutL3_13;

// (* RLOC = "X3Y13" *)
gpc006 gpcL3_13 ({gpcOutL2_8[2],gpcOutL2_9[1],gpcOutL2_10[0],gpcOutL2_40[2],gpcOutL2_41[1],gpcOutL2_42[0]},gpcOutL3_13);
wire [2:0] gpcOutL3_14;

// (* RLOC = "X3Y14" *)
gpc006 gpcL3_14 ({gpcOutL2_9[2],gpcOutL2_10[1],gpcOutL2_11[0],gpcOutL2_41[2],gpcOutL2_42[1],gpcOutL2_43[0]},gpcOutL3_14);
wire [2:0] gpcOutL3_15;

// (* RLOC = "X3Y15" *)
gpc006 gpcL3_15 ({gpcOutL2_10[2],gpcOutL2_11[1],gpcOutL2_12[0],gpcOutL2_42[2],gpcOutL2_43[1],gpcOutL2_44[0]},gpcOutL3_15);
wire [2:0] gpcOutL3_16;

// (* RLOC = "X3Y16" *)
gpc006 gpcL3_16 ({gpcOutL2_11[2],gpcOutL2_12[1],gpcOutL2_18[0],gpcOutL2_43[2],gpcOutL2_44[1],gpcOutL2_60[0]},gpcOutL3_16);
wire [2:0] gpcOutL3_17;

// (* RLOC = "X3Y17" *)
gpc006 gpcL3_17 ({gpcOutL2_25[0],gpcOutL2_33[1],gpcOutL2_52[2],gpcOutL2_77[0],gpcOutL2_87[1],gpcOutL2_116[2]},gpcOutL3_17);
wire [2:0] gpcOutL3_18;

// (* RLOC = "X3Y18" *)
gpc006 gpcL3_18 ({gpcOutL2_19[2],gpcOutL2_26[1],gpcOutL2_27[0],gpcOutL2_63[2],gpcOutL2_78[1],gpcOutL2_79[0]},gpcOutL3_18);
wire [2:0] gpcOutL3_19;

// (* RLOC = "X3Y19" *)
gpc006 gpcL3_19 ({gpcOutL2_13[0],gpcOutL2_16[1],gpcOutL2_27[2],gpcOutL2_53[0],gpcOutL2_58[1],gpcOutL2_79[2]},gpcOutL3_19);
wire [2:0] gpcOutL3_20;

// (* RLOC = "X3Y20" *)
gpc006 gpcL3_20 ({gpcOutL2_7[1],gpcOutL2_14[0],gpcOutL2_17[2],gpcOutL2_39[1],gpcOutL2_54[0],gpcOutL2_59[2]},gpcOutL3_20);
wire [2:0] gpcOutL3_21;

// (* RLOC = "X3Y21" *)
gpc006 gpcL3_21 ({gpcOutL2_18[2],gpcOutL2_20[1],gpcOutL2_21[0],gpcOutL2_60[2],gpcOutL2_64[1],gpcOutL2_65[0]},gpcOutL3_21);
wire [2:0] gpcOutL3_22;

// (* RLOC = "X3Y22" *)
gpc006 gpcL3_22 ({gpcOutL2_20[2],gpcOutL2_21[1],gpcOutL2_22[0],gpcOutL2_64[2],gpcOutL2_65[1],gpcOutL2_66[0]},gpcOutL3_22);
wire [2:0] gpcOutL3_23;

// (* RLOC = "X3Y23" *)
gpc006 gpcL3_23 ({gpcOutL2_21[2],gpcOutL2_22[1],gpcOutL2_23[0],gpcOutL2_65[2],gpcOutL2_66[1],gpcOutL2_67[0]},gpcOutL3_23);
wire [2:0] gpcOutL3_24;

// (* RLOC = "X3Y24" *)
gpc006 gpcL3_24 ({gpcOutL2_22[2],gpcOutL2_23[1],gpcOutL2_24[0],gpcOutL2_66[2],gpcOutL2_67[1],gpcOutL2_68[0]},gpcOutL3_24);
wire [2:0] gpcOutL3_25;

// (* RLOC = "X3Y25" *)
gpc006 gpcL3_25 ({gpcOutL2_23[2],gpcOutL2_24[1],gpcOutL2_37[0],gpcOutL2_67[2],gpcOutL2_68[1],gpcOutL2_91[0]},gpcOutL3_25);
wire [2:0] gpcOutL3_26;

// (* RLOC = "X3Y26" *)
gpc006 gpcL3_26 ({gpcOutL2_25[1],gpcOutL2_33[2],gpcOutL2_34[0],gpcOutL2_77[1],gpcOutL2_87[2],gpcOutL2_88[0]},gpcOutL3_26);
wire [2:0] gpcOutL3_27;

// (* RLOC = "X3Y27" *)
gpc006 gpcL3_27 ({gpcOutL2_19[0],gpcOutL2_25[2],gpcOutL2_34[1],gpcOutL2_63[0],gpcOutL2_77[2],gpcOutL2_88[1]},gpcOutL3_27);
wire [2:0] gpcOutL3_28;

// (* RLOC = "X3Y28" *)
gpc006 gpcL3_28 ({gpcOutL2_19[1],gpcOutL2_26[0],gpcOutL2_34[2],gpcOutL2_63[1],gpcOutL2_78[0],gpcOutL2_88[2]},gpcOutL3_28);
wire [2:0] gpcOutL3_29;

// (* RLOC = "X3Y29" *)
gpc006 gpcL3_29 ({gpcOutL2_16[0],gpcOutL2_26[2],gpcOutL2_27[1],gpcOutL2_58[0],gpcOutL2_78[2],gpcOutL2_79[1]},gpcOutL3_29);
wire [2:0] gpcOutL3_30;

// (* RLOC = "X3Y30" *)
gpc006 gpcL3_30 ({gpcOutL2_49[2],gpcOutL2_61[1],gpcOutL2_69[0],gpcOutL2_105[2],gpcOutL2_127[1],gpcOutL2_137[0]},gpcOutL3_30);
wire [2:0] gpcOutL3_31;

// (* RLOC = "X3Y31" *)
gpc006 gpcL3_31 ({gpcOutL2_50[1],gpcOutL2_56[2],gpcOutL2_57[0],gpcOutL2_114[1],gpcOutL2_122[2],gpcOutL2_123[0]},gpcOutL3_31);
wire [2:0] gpcOutL3_32;

// (* RLOC = "X3Y32" *)
gpc006 gpcL3_32 ({gpcOutL2_38[0],gpcOutL2_50[2],gpcOutL2_57[1],gpcOutL2_94[0],gpcOutL2_114[2],gpcOutL2_123[1]},gpcOutL3_32);
wire [2:0] gpcOutL3_33;

// (* RLOC = "X3Y33" *)
gpc006 gpcL3_33 ({gpcOutL2_38[2],gpcOutL2_51[1],gpcOutL2_52[0],gpcOutL2_94[2],gpcOutL2_115[1],gpcOutL2_116[0]},gpcOutL3_33);
wire [2:0] gpcOutL3_34;

// (* RLOC = "X3Y34" *)
gpc006 gpcL3_34 ({gpcOutL2_33[0],gpcOutL2_51[2],gpcOutL2_52[1],gpcOutL2_87[0],gpcOutL2_115[2],gpcOutL2_116[1]},gpcOutL3_34);
wire [2:0] gpcOutL3_35;

// (* RLOC = "X3Y35" *)
gpc006 gpcL3_35 ({gpcOutL2_24[2],gpcOutL2_37[1],gpcOutL2_45[0],gpcOutL2_68[2],gpcOutL2_91[1],gpcOutL2_101[0]},gpcOutL3_35);
wire [2:0] gpcOutL3_36;

// (* RLOC = "X3Y36" *)
gpc006 gpcL3_36 ({gpcOutL2_37[2],gpcOutL2_45[1],gpcOutL2_46[0],gpcOutL2_91[2],gpcOutL2_101[1],gpcOutL2_102[0]},gpcOutL3_36);
wire [2:0] gpcOutL3_37;

// (* RLOC = "X3Y37" *)
gpc006 gpcL3_37 ({gpcOutL2_45[2],gpcOutL2_46[1],gpcOutL2_47[0],gpcOutL2_101[2],gpcOutL2_102[1],gpcOutL2_103[0]},gpcOutL3_37);
wire [2:0] gpcOutL3_38;

// (* RLOC = "X3Y38" *)
gpc006 gpcL3_38 ({gpcOutL2_46[2],gpcOutL2_47[1],gpcOutL2_48[0],gpcOutL2_102[2],gpcOutL2_103[1],gpcOutL2_104[0]},gpcOutL3_38);
wire [2:0] gpcOutL3_39;

// (* RLOC = "X3Y39" *)
gpc006 gpcL3_39 ({gpcOutL2_47[2],gpcOutL2_48[1],gpcOutL2_49[0],gpcOutL2_103[2],gpcOutL2_104[1],gpcOutL2_105[0]},gpcOutL3_39);
wire [2:0] gpcOutL3_40;

// (* RLOC = "X3Y40" *)
gpc006 gpcL3_40 ({gpcOutL2_48[2],gpcOutL2_49[1],gpcOutL2_61[0],gpcOutL2_104[2],gpcOutL2_105[1],gpcOutL2_127[0]},gpcOutL3_40);
wire [2:0] gpcOutL3_41;

// (* RLOC = "X3Y41" *)
gpc006 gpcL3_41 ({gpcOutL2_74[0],gpcOutL2_85[1],gpcOutL2_113[2],gpcOutL2_150[0],gpcOutL2_163[1],gpcOutL2_201[2]},gpcOutL3_41);
wire [2:0] gpcOutL3_42;

// (* RLOC = "X3Y42" *)
gpc006 gpcL3_42 ({gpcOutL2_62[2],gpcOutL2_75[1],gpcOutL2_76[0],gpcOutL2_130[2],gpcOutL2_151[1],gpcOutL2_152[0]},gpcOutL3_42);
wire [2:0] gpcOutL3_43;

// (* RLOC = "X3Y43" *)
gpc006 gpcL3_43 ({gpcOutL2_50[0],gpcOutL2_56[1],gpcOutL2_76[2],gpcOutL2_114[0],gpcOutL2_122[1],gpcOutL2_152[2]},gpcOutL3_43);
wire [2:0] gpcOutL3_44;

// (* RLOC = "X3Y44" *)
gpc006 gpcL3_44 ({gpcOutL2_38[1],gpcOutL2_51[0],gpcOutL2_57[2],gpcOutL2_94[1],gpcOutL2_115[0],gpcOutL2_123[2]},gpcOutL3_44);
wire [2:0] gpcOutL3_45;

// (* RLOC = "X3Y45" *)
gpc006 gpcL3_45 ({gpcOutL2_81[1],gpcOutL2_82[0],gpcOutL2_90[2],gpcOutL2_157[1],gpcOutL2_158[0],gpcOutL2_168[2]},gpcOutL3_45);
wire [2:0] gpcOutL3_46;

// (* RLOC = "X3Y46" *)
gpc006 gpcL3_46 ({gpcOutL2_61[2],gpcOutL2_69[1],gpcOutL2_70[0],gpcOutL2_127[2],gpcOutL2_137[1],gpcOutL2_138[0]},gpcOutL3_46);
wire [2:0] gpcOutL3_47;

// (* RLOC = "X3Y47" *)
gpc006 gpcL3_47 ({gpcOutL2_69[2],gpcOutL2_70[1],gpcOutL2_71[0],gpcOutL2_137[2],gpcOutL2_138[1],gpcOutL2_139[0]},gpcOutL3_47);
wire [2:0] gpcOutL3_48;

// (* RLOC = "X3Y48" *)
gpc006 gpcL3_48 ({gpcOutL2_70[2],gpcOutL2_71[1],gpcOutL2_72[0],gpcOutL2_138[2],gpcOutL2_139[1],gpcOutL2_140[0]},gpcOutL3_48);
wire [2:0] gpcOutL3_49;

// (* RLOC = "X3Y49" *)
gpc006 gpcL3_49 ({gpcOutL2_71[2],gpcOutL2_72[1],gpcOutL2_73[0],gpcOutL2_139[2],gpcOutL2_140[1],gpcOutL2_141[0]},gpcOutL3_49);
wire [2:0] gpcOutL3_50;

// (* RLOC = "X3Y50" *)
gpc006 gpcL3_50 ({gpcOutL2_72[2],gpcOutL2_73[1],gpcOutL2_92[0],gpcOutL2_140[2],gpcOutL2_141[1],gpcOutL2_170[0]},gpcOutL3_50);
wire [2:0] gpcOutL3_51;

// (* RLOC = "X3Y51" *)
gpc006 gpcL3_51 ({gpcOutL2_74[1],gpcOutL2_85[2],gpcOutL2_86[0],gpcOutL2_150[1],gpcOutL2_163[2],gpcOutL2_164[0]},gpcOutL3_51);
wire [2:0] gpcOutL3_52;

// (* RLOC = "X3Y52" *)
gpc006 gpcL3_52 ({gpcOutL2_62[0],gpcOutL2_74[2],gpcOutL2_86[1],gpcOutL2_130[0],gpcOutL2_150[2],gpcOutL2_164[1]},gpcOutL3_52);
wire [2:0] gpcOutL3_53;

// (* RLOC = "X3Y53" *)
gpc006 gpcL3_53 ({gpcOutL2_62[1],gpcOutL2_75[0],gpcOutL2_86[2],gpcOutL2_130[1],gpcOutL2_151[0],gpcOutL2_164[2]},gpcOutL3_53);
wire [2:0] gpcOutL3_54;

// (* RLOC = "X3Y54" *)
gpc006 gpcL3_54 ({gpcOutL2_56[0],gpcOutL2_75[2],gpcOutL2_76[1],gpcOutL2_122[0],gpcOutL2_151[2],gpcOutL2_152[1]},gpcOutL3_54);
wire [2:0] gpcOutL3_55;

// (* RLOC = "X3Y55" *)
gpc006 gpcL3_55 ({gpcOutL2_80[0],gpcOutL2_89[1],gpcOutL2_119[2],gpcOutL2_156[0],gpcOutL2_167[1],gpcOutL2_207[2]},gpcOutL3_55);
wire [2:0] gpcOutL3_56;

// (* RLOC = "X3Y56" *)
gpc006 gpcL3_56 ({gpcOutL2_80[1],gpcOutL2_89[2],gpcOutL2_90[0],gpcOutL2_156[1],gpcOutL2_167[2],gpcOutL2_168[0]},gpcOutL3_56);
wire [2:0] gpcOutL3_57;

// (* RLOC = "X3Y57" *)
gpc006 gpcL3_57 ({gpcOutL2_80[2],gpcOutL2_81[0],gpcOutL2_90[1],gpcOutL2_156[2],gpcOutL2_157[0],gpcOutL2_168[1]},gpcOutL3_57);
wire [2:0] gpcOutL3_58;

// (* RLOC = "X3Y58" *)
gpc006 gpcL3_58 ({gpcOutL2_81[2],gpcOutL2_82[1],gpcOutL2_83[0],gpcOutL2_157[2],gpcOutL2_158[1],gpcOutL2_159[0]},gpcOutL3_58);
wire [2:0] gpcOutL3_59;

// (* RLOC = "X3Y59" *)
gpc006 gpcL3_59 ({gpcOutL2_82[2],gpcOutL2_83[1],gpcOutL2_84[0],gpcOutL2_158[2],gpcOutL2_159[1],gpcOutL2_160[0]},gpcOutL3_59);
wire [2:0] gpcOutL3_60;

// (* RLOC = "X3Y60" *)
gpc006 gpcL3_60 ({gpcOutL2_83[2],gpcOutL2_84[1],gpcOutL2_96[0],gpcOutL2_159[2],gpcOutL2_160[1],gpcOutL2_176[0]},gpcOutL3_60);
wire [2:0] gpcOutL3_61;

// (* RLOC = "X3Y61" *)
gpc006 gpcL3_61 ({gpcOutL2_100[2],gpcOutL2_126[1],gpcOutL2_132[0],gpcOutL2_180[2],gpcOutL2_216[1],gpcOutL2_224[0]},gpcOutL3_61);
wire [2:0] gpcOutL3_62;

// (* RLOC = "X3Y62" *)
gpc006 gpcL3_62 ({gpcOutL2_110[2],gpcOutL2_128[1],gpcOutL2_142[0],gpcOutL2_190[2],gpcOutL2_218[1],gpcOutL2_234[0]},gpcOutL3_62);
wire [2:0] gpcOutL3_63;

// (* RLOC = "X3Y63" *)
gpc006 gpcL3_63 ({gpcOutL2_111[1],gpcOutL2_120[2],gpcOutL2_121[0],gpcOutL2_199[1],gpcOutL2_210[2],gpcOutL2_211[0]},gpcOutL3_63);
wire [2:0] gpcOutL3_64;

// (* RLOC = "X3Y64" *)
gpc006 gpcL3_64 ({gpcOutL2_93[0],gpcOutL2_111[2],gpcOutL2_121[1],gpcOutL2_173[0],gpcOutL2_199[2],gpcOutL2_211[1]},gpcOutL3_64);
wire [2:0] gpcOutL3_65;

// (* RLOC = "X3Y65" *)
gpc006 gpcL3_65 ({gpcOutL2_93[2],gpcOutL2_112[1],gpcOutL2_113[0],gpcOutL2_173[2],gpcOutL2_200[1],gpcOutL2_201[0]},gpcOutL3_65);
wire [2:0] gpcOutL3_66;

// (* RLOC = "X3Y66" *)
gpc006 gpcL3_66 ({gpcOutL2_85[0],gpcOutL2_112[2],gpcOutL2_113[1],gpcOutL2_163[0],gpcOutL2_200[2],gpcOutL2_201[1]},gpcOutL3_66);
wire [2:0] gpcOutL3_67;

// (* RLOC = "X3Y67" *)
gpc006 gpcL3_67 ({gpcOutL2_117[1],gpcOutL2_124[2],gpcOutL2_125[0],gpcOutL2_205[1],gpcOutL2_214[2],gpcOutL2_215[0]},gpcOutL3_67);
wire [2:0] gpcOutL3_68;

// (* RLOC = "X3Y68" *)
gpc006 gpcL3_68 ({gpcOutL2_95[0],gpcOutL2_117[2],gpcOutL2_125[1],gpcOutL2_175[0],gpcOutL2_205[2],gpcOutL2_215[1]},gpcOutL3_68);
wire [2:0] gpcOutL3_69;

// (* RLOC = "X3Y69" *)
gpc006 gpcL3_69 ({gpcOutL2_95[2],gpcOutL2_118[1],gpcOutL2_119[0],gpcOutL2_175[2],gpcOutL2_206[1],gpcOutL2_207[0]},gpcOutL3_69);
wire [2:0] gpcOutL3_70;

// (* RLOC = "X3Y70" *)
gpc006 gpcL3_70 ({gpcOutL2_89[0],gpcOutL2_118[2],gpcOutL2_119[1],gpcOutL2_167[0],gpcOutL2_206[2],gpcOutL2_207[1]},gpcOutL3_70);
wire [2:0] gpcOutL3_71;

// (* RLOC = "X3Y71" *)
gpc006 gpcL3_71 ({gpcOutL2_84[2],gpcOutL2_96[1],gpcOutL2_97[0],gpcOutL2_160[2],gpcOutL2_176[1],gpcOutL2_177[0]},gpcOutL3_71);
wire [2:0] gpcOutL3_72;

// (* RLOC = "X3Y72" *)
gpc006 gpcL3_72 ({gpcOutL2_96[2],gpcOutL2_97[1],gpcOutL2_98[0],gpcOutL2_176[2],gpcOutL2_177[1],gpcOutL2_178[0]},gpcOutL3_72);
wire [2:0] gpcOutL3_73;

// (* RLOC = "X3Y73" *)
gpc006 gpcL3_73 ({gpcOutL2_97[2],gpcOutL2_98[1],gpcOutL2_99[0],gpcOutL2_177[2],gpcOutL2_178[1],gpcOutL2_179[0]},gpcOutL3_73);
wire [2:0] gpcOutL3_74;

// (* RLOC = "X3Y74" *)
gpc006 gpcL3_74 ({gpcOutL2_98[2],gpcOutL2_99[1],gpcOutL2_100[0],gpcOutL2_178[2],gpcOutL2_179[1],gpcOutL2_180[0]},gpcOutL3_74);
wire [2:0] gpcOutL3_75;

// (* RLOC = "X3Y75" *)
gpc006 gpcL3_75 ({gpcOutL2_99[2],gpcOutL2_100[1],gpcOutL2_126[0],gpcOutL2_179[2],gpcOutL2_180[1],gpcOutL2_216[0]},gpcOutL3_75);
wire [2:0] gpcOutL3_76;

// (* RLOC = "X3Y76" *)
gpc006 gpcL3_76 ({gpcOutL2_73[2],gpcOutL2_92[1],gpcOutL2_106[0],gpcOutL2_141[2],gpcOutL2_170[1],gpcOutL2_186[0]},gpcOutL3_76);
wire [2:0] gpcOutL3_77;

// (* RLOC = "X3Y77" *)
gpc006 gpcL3_77 ({gpcOutL2_92[2],gpcOutL2_106[1],gpcOutL2_107[0],gpcOutL2_170[2],gpcOutL2_186[1],gpcOutL2_187[0]},gpcOutL3_77);
wire [2:0] gpcOutL3_78;

// (* RLOC = "X3Y78" *)
gpc006 gpcL3_78 ({gpcOutL2_106[2],gpcOutL2_107[1],gpcOutL2_108[0],gpcOutL2_186[2],gpcOutL2_187[1],gpcOutL2_188[0]},gpcOutL3_78);
wire [2:0] gpcOutL3_79;

// (* RLOC = "X3Y79" *)
gpc006 gpcL3_79 ({gpcOutL2_107[2],gpcOutL2_108[1],gpcOutL2_109[0],gpcOutL2_187[2],gpcOutL2_188[1],gpcOutL2_189[0]},gpcOutL3_79);
wire [2:0] gpcOutL3_80;

// (* RLOC = "X3Y80" *)
gpc006 gpcL3_80 ({gpcOutL2_108[2],gpcOutL2_109[1],gpcOutL2_110[0],gpcOutL2_188[2],gpcOutL2_189[1],gpcOutL2_190[0]},gpcOutL3_80);
wire [2:0] gpcOutL3_81;

// (* RLOC = "X3Y81" *)
gpc006 gpcL3_81 ({gpcOutL2_109[2],gpcOutL2_110[1],gpcOutL2_128[0],gpcOutL2_189[2],gpcOutL2_190[1],gpcOutL2_218[0]},gpcOutL3_81);
wire [2:0] gpcOutL3_82;

// (* RLOC = "X3Y82" *)
gpc006 gpcL3_82 ({gpcOutL2_147[0],gpcOutL2_161[1],gpcOutL2_198[2],gpcOutL2_247[0],gpcOutL2_263[1],gpcOutL2_318[2]},gpcOutL3_82);
wire [2:0] gpcOutL3_83;

// (* RLOC = "X3Y83" *)
gpc006 gpcL3_83 ({gpcOutL2_129[2],gpcOutL2_148[1],gpcOutL2_149[0],gpcOutL2_221[2],gpcOutL2_248[1],gpcOutL2_249[0]},gpcOutL3_83);
wire [2:0] gpcOutL3_84;

// (* RLOC = "X3Y84" *)
gpc006 gpcL3_84 ({gpcOutL2_111[0],gpcOutL2_120[1],gpcOutL2_149[2],gpcOutL2_199[0],gpcOutL2_210[1],gpcOutL2_249[2]},gpcOutL3_84);
wire [2:0] gpcOutL3_85;

// (* RLOC = "X3Y85" *)
gpc006 gpcL3_85 ({gpcOutL2_93[1],gpcOutL2_112[0],gpcOutL2_121[2],gpcOutL2_173[1],gpcOutL2_200[0],gpcOutL2_211[2]},gpcOutL3_85);
wire [2:0] gpcOutL3_86;

// (* RLOC = "X3Y86" *)
gpc006 gpcL3_86 ({gpcOutL2_153[0],gpcOutL2_165[1],gpcOutL2_204[2],gpcOutL2_253[0],gpcOutL2_267[1],gpcOutL2_322[2]},gpcOutL3_86);
wire [2:0] gpcOutL3_87;

// (* RLOC = "X3Y87" *)
gpc006 gpcL3_87 ({gpcOutL2_131[2],gpcOutL2_154[1],gpcOutL2_155[0],gpcOutL2_223[2],gpcOutL2_254[1],gpcOutL2_255[0]},gpcOutL3_87);
wire [2:0] gpcOutL3_88;

// (* RLOC = "X3Y88" *)
gpc006 gpcL3_88 ({gpcOutL2_117[0],gpcOutL2_124[1],gpcOutL2_155[2],gpcOutL2_205[0],gpcOutL2_214[1],gpcOutL2_255[2]},gpcOutL3_88);
wire [2:0] gpcOutL3_89;

// (* RLOC = "X3Y89" *)
gpc006 gpcL3_89 ({gpcOutL2_95[1],gpcOutL2_118[0],gpcOutL2_125[2],gpcOutL2_175[1],gpcOutL2_206[0],gpcOutL2_215[2]},gpcOutL3_89);
wire [2:0] gpcOutL3_90;

// (* RLOC = "X3Y90" *)
gpc006 gpcL3_90 ({gpcOutL2_126[2],gpcOutL2_132[1],gpcOutL2_133[0],gpcOutL2_216[2],gpcOutL2_224[1],gpcOutL2_225[0]},gpcOutL3_90);
wire [2:0] gpcOutL3_91;

// (* RLOC = "X3Y91" *)
gpc006 gpcL3_91 ({gpcOutL2_132[2],gpcOutL2_133[1],gpcOutL2_134[0],gpcOutL2_224[2],gpcOutL2_225[1],gpcOutL2_226[0]},gpcOutL3_91);
wire [2:0] gpcOutL3_92;

// (* RLOC = "X3Y92" *)
gpc006 gpcL3_92 ({gpcOutL2_133[2],gpcOutL2_134[1],gpcOutL2_135[0],gpcOutL2_225[2],gpcOutL2_226[1],gpcOutL2_227[0]},gpcOutL3_92);
wire [2:0] gpcOutL3_93;

// (* RLOC = "X3Y93" *)
gpc006 gpcL3_93 ({gpcOutL2_134[2],gpcOutL2_135[1],gpcOutL2_136[0],gpcOutL2_226[2],gpcOutL2_227[1],gpcOutL2_228[0]},gpcOutL3_93);
wire [2:0] gpcOutL3_94;

// (* RLOC = "X3Y94" *)
gpc006 gpcL3_94 ({gpcOutL2_135[2],gpcOutL2_136[1],gpcOutL2_169[0],gpcOutL2_227[2],gpcOutL2_228[1],gpcOutL2_271[0]},gpcOutL3_94);
wire [2:0] gpcOutL3_95;

// (* RLOC = "X3Y95" *)
gpc006 gpcL3_95 ({gpcOutL2_128[2],gpcOutL2_142[1],gpcOutL2_143[0],gpcOutL2_218[2],gpcOutL2_234[1],gpcOutL2_235[0]},gpcOutL3_95);
wire [2:0] gpcOutL3_96;

// (* RLOC = "X3Y96" *)
gpc006 gpcL3_96 ({gpcOutL2_142[2],gpcOutL2_143[1],gpcOutL2_144[0],gpcOutL2_234[2],gpcOutL2_235[1],gpcOutL2_236[0]},gpcOutL3_96);
wire [2:0] gpcOutL3_97;

// (* RLOC = "X3Y97" *)
gpc006 gpcL3_97 ({gpcOutL2_143[2],gpcOutL2_144[1],gpcOutL2_145[0],gpcOutL2_235[2],gpcOutL2_236[1],gpcOutL2_237[0]},gpcOutL3_97);
wire [2:0] gpcOutL3_98;

// (* RLOC = "X3Y98" *)
gpc006 gpcL3_98 ({gpcOutL2_144[2],gpcOutL2_145[1],gpcOutL2_146[0],gpcOutL2_236[2],gpcOutL2_237[1],gpcOutL2_238[0]},gpcOutL3_98);
wire [2:0] gpcOutL3_99;

// (* RLOC = "X3Y99" *)
gpc006 gpcL3_99 ({gpcOutL2_145[2],gpcOutL2_146[1],gpcOutL2_171[0],gpcOutL2_237[2],gpcOutL2_238[1],gpcOutL2_273[0]},gpcOutL3_99);
wire [2:0] gpcOutL3_100;

// (* RLOC = "X3Y100" *)
gpc006 gpcL3_100 ({gpcOutL2_147[1],gpcOutL2_161[2],gpcOutL2_162[0],gpcOutL2_247[1],gpcOutL2_263[2],gpcOutL2_264[0]},gpcOutL3_100);
wire [2:0] gpcOutL3_101;

// (* RLOC = "X3Y101" *)
gpc006 gpcL3_101 ({gpcOutL2_129[0],gpcOutL2_147[2],gpcOutL2_162[1],gpcOutL2_221[0],gpcOutL2_247[2],gpcOutL2_264[1]},gpcOutL3_101);
wire [2:0] gpcOutL3_102;

// (* RLOC = "X3Y102" *)
gpc006 gpcL3_102 ({gpcOutL2_129[1],gpcOutL2_148[0],gpcOutL2_162[2],gpcOutL2_221[1],gpcOutL2_248[0],gpcOutL2_264[2]},gpcOutL3_102);
wire [2:0] gpcOutL3_103;

// (* RLOC = "X3Y103" *)
gpc006 gpcL3_103 ({gpcOutL2_120[0],gpcOutL2_148[2],gpcOutL2_149[1],gpcOutL2_210[0],gpcOutL2_248[2],gpcOutL2_249[1]},gpcOutL3_103);
wire [2:0] gpcOutL3_104;

// (* RLOC = "X3Y104" *)
gpc006 gpcL3_104 ({gpcOutL2_153[1],gpcOutL2_165[2],gpcOutL2_166[0],gpcOutL2_253[1],gpcOutL2_267[2],gpcOutL2_268[0]},gpcOutL3_104);
wire [2:0] gpcOutL3_105;

// (* RLOC = "X3Y105" *)
gpc006 gpcL3_105 ({gpcOutL2_131[0],gpcOutL2_153[2],gpcOutL2_166[1],gpcOutL2_223[0],gpcOutL2_253[2],gpcOutL2_268[1]},gpcOutL3_105);
wire [2:0] gpcOutL3_106;

// (* RLOC = "X3Y106" *)
gpc006 gpcL3_106 ({gpcOutL2_131[1],gpcOutL2_154[0],gpcOutL2_166[2],gpcOutL2_223[1],gpcOutL2_254[0],gpcOutL2_268[2]},gpcOutL3_106);
wire [2:0] gpcOutL3_107;

// (* RLOC = "X3Y107" *)
gpc006 gpcL3_107 ({gpcOutL2_124[0],gpcOutL2_154[2],gpcOutL2_155[1],gpcOutL2_214[0],gpcOutL2_254[2],gpcOutL2_255[1]},gpcOutL3_107);
wire [2:0] gpcOutL3_108;

// (* RLOC = "X3Y108" *)
gpc006 gpcL3_108 ({gpcOutL2_185[2],gpcOutL2_217[1],gpcOutL2_229[0],gpcOutL2_289[2],gpcOutL2_326[1],gpcOutL1_603[1]},gpcOutL3_108);
wire [2:0] gpcOutL3_109;

// (* RLOC = "X3Y109" *)
gpc006 gpcL3_109 ({gpcOutL2_195[2],gpcOutL2_219[1],gpcOutL2_239[0],gpcOutL2_299[2],gpcOutL2_328[1],gpcOutL1_607[1]},gpcOutL3_109);
wire [2:0] gpcOutL3_110;

// (* RLOC = "X3Y110" *)
gpc006 gpcL3_110 ({gpcOutL2_196[1],gpcOutL2_208[2],gpcOutL2_209[0],gpcOutL2_307[1],gpcOutL2_317[3],gpcOutL2_333[0]},gpcOutL3_110);
wire [2:0] gpcOutL3_111;

// (* RLOC = "X3Y111" *)
gpc006 gpcL3_111 ({gpcOutL2_172[0],gpcOutL2_196[2],gpcOutL2_209[1],gpcOutL2_276[0],gpcOutL2_307[2],gpcOutL2_333[1]},gpcOutL3_111);
wire [2:0] gpcOutL3_112;

// (* RLOC = "X3Y112" *)
gpc006 gpcL3_112 ({gpcOutL2_172[2],gpcOutL2_197[1],gpcOutL2_198[0],gpcOutL2_276[2],gpcOutL2_308[1],gpcOutL2_318[0]},gpcOutL3_112);
wire [2:0] gpcOutL3_113;

// (* RLOC = "X3Y113" *)
gpc006 gpcL3_113 ({gpcOutL2_161[0],gpcOutL2_197[2],gpcOutL2_198[1],gpcOutL2_263[0],gpcOutL2_308[2],gpcOutL2_318[1]},gpcOutL3_113);
wire [2:0] gpcOutL3_114;

// (* RLOC = "X3Y114" *)
gpc006 gpcL3_114 ({gpcOutL2_202[1],gpcOutL2_212[2],gpcOutL2_213[0],gpcOutL2_311[1],gpcOutL2_321[3],gpcOutL2_337[0]},gpcOutL3_114);
wire [2:0] gpcOutL3_115;

// (* RLOC = "X3Y115" *)
gpc006 gpcL3_115 ({gpcOutL2_174[0],gpcOutL2_202[2],gpcOutL2_213[1],gpcOutL2_278[0],gpcOutL2_311[2],gpcOutL2_337[1]},gpcOutL3_115);
wire [2:0] gpcOutL3_116;

// (* RLOC = "X3Y116" *)
gpc006 gpcL3_116 ({gpcOutL2_174[2],gpcOutL2_203[1],gpcOutL2_204[0],gpcOutL2_278[2],gpcOutL2_312[1],gpcOutL2_322[0]},gpcOutL3_116);
wire [2:0] gpcOutL3_117;

// (* RLOC = "X3Y117" *)
gpc006 gpcL3_117 ({gpcOutL2_165[0],gpcOutL2_203[2],gpcOutL2_204[1],gpcOutL2_267[0],gpcOutL2_312[2],gpcOutL2_322[1]},gpcOutL3_117);
wire [2:0] gpcOutL3_118;

// (* RLOC = "X3Y118" *)
gpc006 gpcL3_118 ({gpcOutL2_136[2],gpcOutL2_169[1],gpcOutL2_181[0],gpcOutL2_228[2],gpcOutL2_271[1],gpcOutL2_285[0]},gpcOutL3_118);
wire [2:0] gpcOutL3_119;

// (* RLOC = "X3Y119" *)
gpc006 gpcL3_119 ({gpcOutL2_169[2],gpcOutL2_181[1],gpcOutL2_182[0],gpcOutL2_271[2],gpcOutL2_285[1],gpcOutL2_286[0]},gpcOutL3_119);
wire [2:0] gpcOutL3_120;

// (* RLOC = "X3Y120" *)
gpc006 gpcL3_120 ({gpcOutL2_181[2],gpcOutL2_182[1],gpcOutL2_183[0],gpcOutL2_285[2],gpcOutL2_286[1],gpcOutL2_287[0]},gpcOutL3_120);
wire [2:0] gpcOutL3_121;

// (* RLOC = "X3Y121" *)
gpc006 gpcL3_121 ({gpcOutL2_182[2],gpcOutL2_183[1],gpcOutL2_184[0],gpcOutL2_286[2],gpcOutL2_287[1],gpcOutL2_288[0]},gpcOutL3_121);
wire [2:0] gpcOutL3_122;

// (* RLOC = "X3Y122" *)
gpc006 gpcL3_122 ({gpcOutL2_183[2],gpcOutL2_184[1],gpcOutL2_185[0],gpcOutL2_287[2],gpcOutL2_288[1],gpcOutL2_289[0]},gpcOutL3_122);
wire [2:0] gpcOutL3_123;

// (* RLOC = "X3Y123" *)
gpc006 gpcL3_123 ({gpcOutL2_184[2],gpcOutL2_185[1],gpcOutL2_217[0],gpcOutL2_288[2],gpcOutL2_289[1],gpcOutL2_326[0]},gpcOutL3_123);
wire [2:0] gpcOutL3_124;

// (* RLOC = "X3Y124" *)
gpc006 gpcL3_124 ({gpcOutL2_146[2],gpcOutL2_171[1],gpcOutL2_191[0],gpcOutL2_238[2],gpcOutL2_273[1],gpcOutL2_295[0]},gpcOutL3_124);
wire [2:0] gpcOutL3_125;

// (* RLOC = "X3Y125" *)
gpc006 gpcL3_125 ({gpcOutL2_171[2],gpcOutL2_191[1],gpcOutL2_192[0],gpcOutL2_273[2],gpcOutL2_295[1],gpcOutL2_296[0]},gpcOutL3_125);
wire [2:0] gpcOutL3_126;

// (* RLOC = "X3Y126" *)
gpc006 gpcL3_126 ({gpcOutL2_191[2],gpcOutL2_192[1],gpcOutL2_193[0],gpcOutL2_295[2],gpcOutL2_296[1],gpcOutL2_297[0]},gpcOutL3_126);
wire [2:0] gpcOutL3_127;

// (* RLOC = "X3Y127" *)
gpc006 gpcL3_127 ({gpcOutL2_192[2],gpcOutL2_193[1],gpcOutL2_194[0],gpcOutL2_296[2],gpcOutL2_297[1],gpcOutL2_298[0]},gpcOutL3_127);
wire [2:0] gpcOutL3_128;

// (* RLOC = "X3Y128" *)
gpc006 gpcL3_128 ({gpcOutL2_193[2],gpcOutL2_194[1],gpcOutL2_195[0],gpcOutL2_297[2],gpcOutL2_298[1],gpcOutL2_299[0]},gpcOutL3_128);
wire [2:0] gpcOutL3_129;

// (* RLOC = "X3Y129" *)
gpc006 gpcL3_129 ({gpcOutL2_194[2],gpcOutL2_195[1],gpcOutL2_219[0],gpcOutL2_298[2],gpcOutL2_299[1],gpcOutL2_328[0]},gpcOutL3_129);
wire [2:0] gpcOutL3_130;

// (* RLOC = "X3Y130" *)
gpc015 gpcL3_130 ({gpcOutL2_244[1],gpcOutL2_244[0],gpcOutL2_261[1],gpcOutL2_316[2],pp12[1],pp13[0]},gpcOutL3_130);
wire [2:0] gpcOutL3_131;

// (* RLOC = "X3Y131" *)
gpc015 gpcL3_131 ({gpcOutL2_208[0],gpcOutL2_220[2],gpcOutL2_245[1],gpcOutL2_246[0],gpcOutL2_317[0],gpcOutL2_332[2]},gpcOutL3_131);
wire [2:0] gpcOutL3_132;

// (* RLOC = "X3Y132" *)
gpc005 gpcL3_132 ({gpcOutL2_196[0],gpcOutL2_208[1],gpcOutL2_246[2],gpcOutL2_307[0],gpcOutL2_317[2]},gpcOutL3_132);
wire [2:0] gpcOutL3_133;

// (* RLOC = "X3Y133" *)
gpc005 gpcL3_133 ({gpcOutL2_172[1],gpcOutL2_197[0],gpcOutL2_209[2],gpcOutL2_276[1],gpcOutL2_308[0]},gpcOutL3_133);
wire [2:0] gpcOutL3_134;

// (* RLOC = "X3Y134" *)
gpc015 gpcL3_134 ({gpcOutL2_250[1],gpcOutL2_250[0],gpcOutL2_265[1],gpcOutL2_320[2],pp36[1],pp37[0]},gpcOutL3_134);
wire [2:0] gpcOutL3_135;

// (* RLOC = "X3Y135" *)
gpc015 gpcL3_135 ({gpcOutL2_212[0],gpcOutL2_222[2],gpcOutL2_251[1],gpcOutL2_252[0],gpcOutL2_321[0],gpcOutL2_336[2]},gpcOutL3_135);
wire [2:0] gpcOutL3_136;

// (* RLOC = "X3Y136" *)
gpc005 gpcL3_136 ({gpcOutL2_202[0],gpcOutL2_212[1],gpcOutL2_252[2],gpcOutL2_311[0],gpcOutL2_321[2]},gpcOutL3_136);
wire [2:0] gpcOutL3_137;

// (* RLOC = "X3Y137" *)
gpc005 gpcL3_137 ({gpcOutL2_174[1],gpcOutL2_203[0],gpcOutL2_213[2],gpcOutL2_278[1],gpcOutL2_312[0]},gpcOutL3_137);
wire [2:0] gpcOutL3_138;

// (* RLOC = "X3Y138" *)
gpc015 gpcL3_138 ({gpcOutL2_257[2],gpcOutL2_257[1],gpcOutL2_258[0],gpcOutL2_270[2],gpcOutL2_350[3],gpcOutL2_351[0]},gpcOutL3_138);
wire [2:0] gpcOutL3_139;

// (* RLOC = "X3Y139" *)
gpc015 gpcL3_139 ({gpcOutL2_229[2],gpcOutL2_217[2],gpcOutL2_229[1],gpcOutL2_230[0],gpcOutL2_326[2],gpcOutL2_342[0]},gpcOutL3_139);
wire [2:0] gpcOutL3_140;

// (* RLOC = "X3Y140" *)
gpc015 gpcL3_140 ({gpcOutL2_231[2],gpcOutL2_230[2],gpcOutL2_231[1],gpcOutL2_232[0],gpcOutL2_342[2],gpcOutL2_343[0]},gpcOutL3_140);
wire [2:0] gpcOutL3_141;

// (* RLOC = "X3Y141" *)
gpc015 gpcL3_141 ({gpcOutL2_233[2],gpcOutL2_232[2],gpcOutL2_233[1],gpcOutL2_272[0],gpcOutL2_343[2],pp63[27]},gpcOutL3_141);
wire [2:0] gpcOutL3_142;

// (* RLOC = "X3Y142" *)
gpc015 gpcL3_142 ({gpcOutL2_239[2],gpcOutL2_219[2],gpcOutL2_239[1],gpcOutL2_240[0],gpcOutL2_328[2],gpcOutL2_346[0]},gpcOutL3_142);
wire [2:0] gpcOutL3_143;

// (* RLOC = "X3Y143" *)
gpc015 gpcL3_143 ({gpcOutL2_241[2],gpcOutL2_240[2],gpcOutL2_241[1],gpcOutL2_242[0],gpcOutL2_346[2],gpcOutL2_347[0]},gpcOutL3_143);
wire [2:0] gpcOutL3_144;

// (* RLOC = "X3Y144" *)
gpc015 gpcL3_144 ({gpcOutL2_243[2],gpcOutL2_242[2],gpcOutL2_243[1],gpcOutL2_274[0],gpcOutL2_347[2],pp63[51]},gpcOutL3_144);
wire [2:0] gpcOutL3_145;

// (* RLOC = "X3Y145" *)
gpc014 gpcL3_145 ({gpcOutL2_220[1],gpcOutL2_220[0],gpcOutL2_244[2],gpcOutL2_262[1],gpcOutL2_332[0]},gpcOutL3_145);
wire [2:0] gpcOutL3_146;

// (* RLOC = "X3Y146" *)
gpc014 gpcL3_146 ({gpcOutL2_222[1],gpcOutL2_222[0],gpcOutL2_250[2],gpcOutL2_266[1],gpcOutL2_336[0]},gpcOutL3_146);
wire [2:0] gpcOutL3_147;

// (* RLOC = "X3Y147" *)
gpc014 gpcL3_147 ({gpcOutL2_256[1],gpcOutL2_256[0],gpcOutL2_269[1],gpcOutL2_324[2],gpcOutL2_350[0]},gpcOutL3_147);
wire [2:0] gpcOutL3_148;

// (* RLOC = "X3Y148" *)
gpc023 gpcL3_148 ({gpcOutL2_256[2],gpcOutL2_257[0],gpcOutL2_269[2],gpcOutL2_270[0],gpcOutL2_350[1]},gpcOutL3_148);
wire [2:0] gpcOutL3_149;

// (* RLOC = "X3Y149" *)
gpc014 gpcL3_149 ({gpcOutL2_259[2],gpcOutL2_258[2],gpcOutL2_259[1],gpcOutL2_260[0],gpcOutL2_351[2]},gpcOutL3_149);
wire [2:0] gpcOutL3_150;

// (* RLOC = "X3Y150" *)
gpc014 gpcL3_150 ({gpcOutL2_325[2],gpcOutL2_284[2],gpcOutL2_325[1],gpcOutL1_601[1],gpcOutL1_621[0]},gpcOutL3_150);
wire [1:0] gpcOutL3_151;

// (* RLOC = "X3Y151" *)
gpc003 gpcL3_151 ({gpcOutL2_230[1],gpcOutL2_231[0],gpcOutL2_342[1]},gpcOutL3_151);
wire [1:0] gpcOutL3_152;

// (* RLOC = "X3Y152" *)
gpc003 gpcL3_152 ({gpcOutL2_232[1],gpcOutL2_233[0],gpcOutL2_343[1]},gpcOutL3_152);
wire [2:0] gpcOutL3_153;

// (* RLOC = "X3Y153" *)
gpc014 gpcL3_153 ({gpcOutL2_327[2],gpcOutL2_294[2],gpcOutL2_327[1],gpcOutL1_605[1],gpcOutL1_625[0]},gpcOutL3_153);
wire [1:0] gpcOutL3_154;

// (* RLOC = "X3Y154" *)
gpc003 gpcL3_154 ({gpcOutL2_240[1],gpcOutL2_241[0],gpcOutL2_346[1]},gpcOutL3_154);
wire [1:0] gpcOutL3_155;

// (* RLOC = "X3Y155" *)
gpc003 gpcL3_155 ({gpcOutL2_242[1],gpcOutL2_243[0],gpcOutL2_347[1]},gpcOutL3_155);
wire [2:0] gpcOutL3_156;

// (* RLOC = "X3Y156" *)
gpc014 gpcL3_156 ({gpcOutL2_329[2],gpcOutL2_304[2],gpcOutL2_329[1],gpcOutL1_609[1],gpcOutL1_629[0]},gpcOutL3_156);
wire [2:0] gpcOutL3_157;

// (* RLOC = "X3Y157" *)
gpc023 gpcL3_157 ({gpcOutL2_275[0],gpcOutL2_305[2],gpcOutL2_305[1],gpcOutL2_315[3],gpcOutL2_331[0]},gpcOutL3_157);
wire [2:0] gpcOutL3_158;

// (* RLOC = "X3Y158" *)
gpc023 gpcL3_158 ({gpcOutL2_261[0],gpcOutL2_306[2],gpcOutL2_275[2],gpcOutL2_306[1],gpcOutL2_316[0]},gpcOutL3_158);
wire [1:0] gpcOutL3_159;

// (* RLOC = "X3Y159" *)
gpc003 gpcL3_159 ({gpcOutL2_261[2],gpcOutL2_262[0],gpcOutL1_652[0]},gpcOutL3_159);
wire [1:0] gpcOutL3_160;

// (* RLOC = "X3Y160" *)
gpc003 gpcL3_160 ({gpcOutL2_245[0],gpcOutL2_262[2],gpcOutL2_332[1]},gpcOutL3_160);
wire [1:0] gpcOutL3_161;

// (* RLOC = "X3Y161" *)
gpc003 gpcL3_161 ({gpcOutL2_245[2],gpcOutL2_246[1],gpcOutL2_317[1]},gpcOutL3_161);
wire [2:0] gpcOutL3_162;

// (* RLOC = "X3Y162" *)
gpc023 gpcL3_162 ({gpcOutL2_277[0],gpcOutL2_309[2],gpcOutL2_309[1],gpcOutL2_319[3],gpcOutL2_335[0]},gpcOutL3_162);
wire [2:0] gpcOutL3_163;

// (* RLOC = "X3Y163" *)
gpc023 gpcL3_163 ({gpcOutL2_265[0],gpcOutL2_310[2],gpcOutL2_277[2],gpcOutL2_310[1],gpcOutL2_320[0]},gpcOutL3_163);
wire [1:0] gpcOutL3_164;

// (* RLOC = "X3Y164" *)
gpc003 gpcL3_164 ({gpcOutL2_265[2],gpcOutL2_266[0],gpcOutL1_656[0]},gpcOutL3_164);
wire [1:0] gpcOutL3_165;

// (* RLOC = "X3Y165" *)
gpc003 gpcL3_165 ({gpcOutL2_251[0],gpcOutL2_266[2],gpcOutL2_336[1]},gpcOutL3_165);
wire [1:0] gpcOutL3_166;

// (* RLOC = "X3Y166" *)
gpc003 gpcL3_166 ({gpcOutL2_251[2],gpcOutL2_252[1],gpcOutL2_321[1]},gpcOutL3_166);
wire [2:0] gpcOutL3_167;

// (* RLOC = "X3Y167" *)
gpc023 gpcL3_167 ({gpcOutL2_279[0],gpcOutL2_313[2],gpcOutL2_313[1],gpcOutL2_323[3],gpcOutL2_339[0]},gpcOutL3_167);
wire [2:0] gpcOutL3_168;

// (* RLOC = "X3Y168" *)
gpc023 gpcL3_168 ({gpcOutL2_269[0],gpcOutL2_314[2],gpcOutL2_279[2],gpcOutL2_314[1],gpcOutL2_324[0]},gpcOutL3_168);
wire [1:0] gpcOutL3_169;

// (* RLOC = "X3Y169" *)
gpc003 gpcL3_169 ({gpcOutL2_258[1],gpcOutL2_259[0],gpcOutL2_351[1]},gpcOutL3_169);
wire [2:0] gpcOutL3_170;

// (* RLOC = "X3Y170" *)
gpc023 gpcL3_170 ({gpcOutL2_260[2],gpcOutL2_280[1],gpcOutL2_260[1],gpcOutL2_280[0],gpcOutL2_351[3]},gpcOutL3_170);
wire [2:0] gpcOutL3_171;

// (* RLOC = "X3Y171" *)
gpc023 gpcL3_171 ({gpcOutL2_281[2],gpcOutL2_282[1],gpcOutL2_280[2],gpcOutL2_281[1],gpcOutL2_282[0]},gpcOutL3_171);
wire [2:0] gpcOutL3_172;

// (* RLOC = "X3Y172" *)
gpc023 gpcL3_172 ({gpcOutL2_283[2],gpcOutL2_284[1],gpcOutL2_282[2],gpcOutL2_283[1],gpcOutL2_284[0]},gpcOutL3_172);
wire [2:0] gpcOutL3_173;

// (* RLOC = "X3Y173" *)
gpc023 gpcL3_173 ({gpcOutL2_290[2],gpcOutL2_291[1],gpcOutL2_272[2],gpcOutL2_290[1],gpcOutL2_291[0]},gpcOutL3_173);
wire [2:0] gpcOutL3_174;

// (* RLOC = "X3Y174" *)
gpc023 gpcL3_174 ({gpcOutL2_292[2],gpcOutL2_293[1],gpcOutL2_291[2],gpcOutL2_292[1],gpcOutL2_293[0]},gpcOutL3_174);
wire [1:0] gpcOutL3_175;

// (* RLOC = "X3Y175" *)
gpc003 gpcL3_175 ({gpcOutL2_293[2],gpcOutL2_294[1],gpcOutL2_327[0]},gpcOutL3_175);
wire [2:0] gpcOutL3_176;

// (* RLOC = "X3Y176" *)
gpc023 gpcL3_176 ({gpcOutL2_300[2],gpcOutL2_301[1],gpcOutL2_274[2],gpcOutL2_300[1],gpcOutL2_301[0]},gpcOutL3_176);
wire [2:0] gpcOutL3_177;

// (* RLOC = "X3Y177" *)
gpc023 gpcL3_177 ({gpcOutL2_302[2],gpcOutL2_303[1],gpcOutL2_301[2],gpcOutL2_302[1],gpcOutL2_303[0]},gpcOutL3_177);
wire [1:0] gpcOutL3_178;

// (* RLOC = "X3Y178" *)
gpc003 gpcL3_178 ({gpcOutL2_303[2],gpcOutL2_304[1],gpcOutL2_329[0]},gpcOutL3_178);
wire [3:0] gpcOutL3_179;

// (* RLOC = "X3Y179" *)
gpc212 gpcL3_179 ({gpcOutL2_305[0],gpcOutL2_315[2],gpcOutL2_315[1],gpcOutL2_315[0],gpcOutL2_330[2]},gpcOutL3_179);
wire [3:0] gpcOutL3_180;

// (* RLOC = "X3Y180" *)
gpc212 gpcL3_180 ({gpcOutL2_309[0],gpcOutL2_319[2],gpcOutL2_319[1],gpcOutL2_319[0],gpcOutL2_334[2]},gpcOutL3_180);
wire [3:0] gpcOutL3_181;

// (* RLOC = "X3Y181" *)
gpc212 gpcL3_181 ({gpcOutL2_313[0],gpcOutL2_323[2],gpcOutL2_323[1],gpcOutL2_323[0],gpcOutL2_338[2]},gpcOutL3_181);
wire [3:0] gpcOutL3_182;

// (* RLOC = "X3Y182" *)
gpc222 gpcL3_182 ({gpcOutL2_341[1],pp63[14],gpcOutL2_340[2],gpcOutL2_341[0],gpcOutL2_340[1],gpcOutL1_663[0]},gpcOutL3_182);
wire [3:0] gpcOutL3_183;

// (* RLOC = "X3Y183" *)
gpc222 gpcL3_183 ({gpcOutL2_345[1],pp63[38],gpcOutL2_344[2],gpcOutL2_345[0],gpcOutL2_344[1],gpcOutL1_667[0]},gpcOutL3_183);
wire [3:0] gpcOutL3_184;

// (* RLOC = "X3Y184" *)
gpc222 gpcL3_184 ({gpcOutL2_349[1],pp63[62],gpcOutL2_348[2],gpcOutL2_349[0],gpcOutL2_348[1],gpcOutL1_671[0]},gpcOutL3_184);
wire [2:0] gpcOutL4_0;

// (* RLOC = "X4Y0" *)
gpc006 gpcL4_0 ({gpcOutL3_1[2],gpcOutL3_2[1],gpcOutL3_3[0],gpcOutL3_55[2],gpcOutL3_56[1],gpcOutL3_57[0]},gpcOutL4_0);
wire [2:0] gpcOutL4_1;

// (* RLOC = "X4Y1" *)
gpc006 gpcL4_1 ({gpcOutL3_8[2],gpcOutL3_9[1],gpcOutL3_20[0],gpcOutL3_67[2],gpcOutL3_68[1],gpcOutL3_89[0]},gpcOutL4_1);
wire [2:0] gpcOutL4_2;

// (* RLOC = "X4Y2" *)
gpc006 gpcL4_2 ({gpcOutL3_0[2],gpcOutL3_4[1],gpcOutL3_5[0],gpcOutL3_45[2],gpcOutL3_58[1],gpcOutL3_59[0]},gpcOutL4_2);
wire [2:0] gpcOutL4_3;

// (* RLOC = "X4Y3" *)
gpc006 gpcL4_3 ({gpcOutL3_5[2],gpcOutL3_6[1],gpcOutL3_12[0],gpcOutL3_59[2],gpcOutL3_60[1],gpcOutL3_71[0]},gpcOutL4_3);
wire [2:0] gpcOutL4_4;

// (* RLOC = "X4Y4" *)
gpc006 gpcL4_4 ({gpcOutL3_23[2],gpcOutL3_24[1],gpcOutL3_25[0],gpcOutL3_92[2],gpcOutL3_93[1],gpcOutL3_94[0]},gpcOutL4_4);
wire [2:0] gpcOutL4_5;

// (* RLOC = "X4Y5" *)
gpc006 gpcL4_5 ({gpcOutL3_17[0],gpcOutL3_33[2],gpcOutL3_34[1],gpcOutL3_86[0],gpcOutL3_116[2],gpcOutL3_117[1]},gpcOutL4_5);
wire [2:0] gpcOutL4_6;

// (* RLOC = "X4Y6" *)
gpc006 gpcL4_6 ({gpcOutL3_8[0],gpcOutL3_19[1],gpcOutL3_29[2],gpcOutL3_67[0],gpcOutL3_88[1],gpcOutL3_107[2]},gpcOutL4_6);
wire [2:0] gpcOutL4_7;

// (* RLOC = "X4Y7" *)
gpc006 gpcL4_7 ({gpcOutL3_8[1],gpcOutL3_9[0],gpcOutL3_19[2],gpcOutL3_67[1],gpcOutL3_68[0],gpcOutL3_88[2]},gpcOutL4_7);
wire [2:0] gpcOutL4_8;

// (* RLOC = "X4Y8" *)
gpc006 gpcL4_8 ({gpcOutL3_10[1],gpcOutL3_11[0],gpcOutL3_20[2],gpcOutL3_69[1],gpcOutL3_70[0],gpcOutL3_89[2]},gpcOutL4_8);
wire [2:0] gpcOutL4_9;

// (* RLOC = "X4Y9" *)
gpc006 gpcL4_9 ({gpcOutL3_1[0],gpcOutL3_10[2],gpcOutL3_11[1],gpcOutL3_55[0],gpcOutL3_69[2],gpcOutL3_70[1]},gpcOutL4_9);
wire [2:0] gpcOutL4_10;

// (* RLOC = "X4Y10" *)
gpc006 gpcL4_10 ({gpcOutL3_1[1],gpcOutL3_2[0],gpcOutL3_11[2],gpcOutL3_55[1],gpcOutL3_56[0],gpcOutL3_70[2]},gpcOutL4_10);
wire [2:0] gpcOutL4_11;

// (* RLOC = "X4Y11" *)
gpc006 gpcL4_11 ({gpcOutL3_0[0],gpcOutL3_2[2],gpcOutL3_3[1],gpcOutL3_45[0],gpcOutL3_56[2],gpcOutL3_57[1]},gpcOutL4_11);
wire [2:0] gpcOutL4_12;

// (* RLOC = "X4Y12" *)
gpc006 gpcL4_12 ({gpcOutL3_0[1],gpcOutL3_3[2],gpcOutL3_4[0],gpcOutL3_45[1],gpcOutL3_57[2],gpcOutL3_58[0]},gpcOutL4_12);
wire [2:0] gpcOutL4_13;

// (* RLOC = "X4Y13" *)
gpc006 gpcL4_13 ({gpcOutL3_4[2],gpcOutL3_5[1],gpcOutL3_6[0],gpcOutL3_58[2],gpcOutL3_59[1],gpcOutL3_60[0]},gpcOutL4_13);
wire [2:0] gpcOutL4_14;

// (* RLOC = "X4Y14" *)
gpc006 gpcL4_14 ({gpcOutL3_6[2],gpcOutL3_12[1],gpcOutL3_13[0],gpcOutL3_60[2],gpcOutL3_71[1],gpcOutL3_72[0]},gpcOutL4_14);
wire [2:0] gpcOutL4_15;

// (* RLOC = "X4Y15" *)
gpc006 gpcL4_15 ({gpcOutL3_12[2],gpcOutL3_13[1],gpcOutL3_14[0],gpcOutL3_71[2],gpcOutL3_72[1],gpcOutL3_73[0]},gpcOutL4_15);
wire [2:0] gpcOutL4_16;

// (* RLOC = "X4Y16" *)
gpc006 gpcL4_16 ({gpcOutL3_13[2],gpcOutL3_14[1],gpcOutL3_15[0],gpcOutL3_72[2],gpcOutL3_73[1],gpcOutL3_74[0]},gpcOutL4_16);
wire [2:0] gpcOutL4_17;

// (* RLOC = "X4Y17" *)
gpc006 gpcL4_17 ({gpcOutL3_14[2],gpcOutL3_15[1],gpcOutL3_16[0],gpcOutL3_73[2],gpcOutL3_74[1],gpcOutL3_75[0]},gpcOutL4_17);
wire [2:0] gpcOutL4_18;

// (* RLOC = "X4Y18" *)
gpc006 gpcL4_18 ({gpcOutL3_7[0],gpcOutL3_15[2],gpcOutL3_16[1],gpcOutL3_61[0],gpcOutL3_74[2],gpcOutL3_75[1]},gpcOutL4_18);
wire [2:0] gpcOutL4_19;

// (* RLOC = "X4Y19" *)
gpc006 gpcL4_19 ({gpcOutL3_7[1],gpcOutL3_16[2],gpcOutL3_21[0],gpcOutL3_61[1],gpcOutL3_75[2],gpcOutL3_90[0]},gpcOutL4_19);
wire [2:0] gpcOutL4_20;

// (* RLOC = "X4Y20" *)
gpc006 gpcL4_20 ({gpcOutL3_7[2],gpcOutL3_21[1],gpcOutL3_22[0],gpcOutL3_61[2],gpcOutL3_90[1],gpcOutL3_91[0]},gpcOutL4_20);
wire [2:0] gpcOutL4_21;

// (* RLOC = "X4Y21" *)
gpc006 gpcL4_21 ({gpcOutL3_17[1],gpcOutL3_26[0],gpcOutL3_34[2],gpcOutL3_86[1],gpcOutL3_104[0],gpcOutL3_117[2]},gpcOutL4_21);
wire [2:0] gpcOutL4_22;

// (* RLOC = "X4Y22" *)
gpc006 gpcL4_22 ({gpcOutL3_17[2],gpcOutL3_26[1],gpcOutL3_27[0],gpcOutL3_86[2],gpcOutL3_104[1],gpcOutL3_105[0]},gpcOutL4_22);
wire [2:0] gpcOutL4_23;

// (* RLOC = "X4Y23" *)
gpc006 gpcL4_23 ({gpcOutL3_26[2],gpcOutL3_27[1],gpcOutL3_28[0],gpcOutL3_104[2],gpcOutL3_105[1],gpcOutL3_106[0]},gpcOutL4_23);
wire [2:0] gpcOutL4_24;

// (* RLOC = "X4Y24" *)
gpc006 gpcL4_24 ({gpcOutL3_18[0],gpcOutL3_27[2],gpcOutL3_28[1],gpcOutL3_87[0],gpcOutL3_105[2],gpcOutL3_106[1]},gpcOutL4_24);
wire [2:0] gpcOutL4_25;

// (* RLOC = "X4Y25" *)
gpc006 gpcL4_25 ({gpcOutL3_18[1],gpcOutL3_28[2],gpcOutL3_29[0],gpcOutL3_87[1],gpcOutL3_106[2],gpcOutL3_107[0]},gpcOutL4_25);
wire [2:0] gpcOutL4_26;

// (* RLOC = "X4Y26" *)
gpc006 gpcL4_26 ({gpcOutL3_18[2],gpcOutL3_19[0],gpcOutL3_29[1],gpcOutL3_87[2],gpcOutL3_88[0],gpcOutL3_107[1]},gpcOutL4_26);
wire [2:0] gpcOutL4_27;

// (* RLOC = "X4Y27" *)
gpc006 gpcL4_27 ({gpcOutL3_9[2],gpcOutL3_10[0],gpcOutL3_20[1],gpcOutL3_68[2],gpcOutL3_69[0],gpcOutL3_89[1]},gpcOutL4_27);
wire [2:0] gpcOutL4_28;

// (* RLOC = "X4Y28" *)
gpc006 gpcL4_28 ({gpcOutL3_21[2],gpcOutL3_22[1],gpcOutL3_23[0],gpcOutL3_90[2],gpcOutL3_91[1],gpcOutL3_92[0]},gpcOutL4_28);
wire [2:0] gpcOutL4_29;

// (* RLOC = "X4Y29" *)
gpc006 gpcL4_29 ({gpcOutL3_22[2],gpcOutL3_23[1],gpcOutL3_24[0],gpcOutL3_91[2],gpcOutL3_92[1],gpcOutL3_93[0]},gpcOutL4_29);
wire [2:0] gpcOutL4_30;

// (* RLOC = "X4Y30" *)
gpc006 gpcL4_30 ({gpcOutL3_30[0],gpcOutL3_39[2],gpcOutL3_40[1],gpcOutL3_108[0],gpcOutL3_122[2],gpcOutL3_123[1]},gpcOutL4_30);
wire [2:0] gpcOutL4_31;

// (* RLOC = "X4Y31" *)
gpc006 gpcL4_31 ({gpcOutL3_30[2],gpcOutL3_46[1],gpcOutL3_47[0],gpcOutL3_108[2],gpcOutL3_139[1],gpcOutL3_151[0]},gpcOutL4_31);
wire [2:0] gpcOutL4_32;

// (* RLOC = "X4Y32" *)
gpc006 gpcL4_32 ({gpcOutL3_63[2],gpcOutL3_64[1],gpcOutL3_85[0],gpcOutL3_162[2],gpcOutL2_277[1],gpcOutL2_310[0]},gpcOutL4_32);
wire [2:0] gpcOutL4_33;

// (* RLOC = "X4Y33" *)
gpc006 gpcL4_33 ({gpcOutL3_41[2],gpcOutL3_51[1],gpcOutL3_52[0],gpcOutL3_134[2],gpcOutL3_146[0],gpcOutL3_164[1]},gpcOutL4_33);
wire [2:0] gpcOutL4_34;

// (* RLOC = "X4Y34" *)
gpc006 gpcL4_34 ({gpcOutL3_42[0],gpcOutL3_52[2],gpcOutL3_53[1],gpcOutL3_135[0],gpcOutL3_146[2],gpcOutL3_165[1]},gpcOutL4_34);
wire [2:0] gpcOutL4_35;

// (* RLOC = "X4Y35" *)
gpc006 gpcL4_35 ({gpcOutL3_42[2],gpcOutL3_43[0],gpcOutL3_54[1],gpcOutL3_135[2],gpcOutL3_136[0],gpcOutL3_166[1]},gpcOutL4_35);
wire [2:0] gpcOutL4_36;

// (* RLOC = "X4Y36" *)
gpc006 gpcL4_36 ({gpcOutL3_31[1],gpcOutL3_32[0],gpcOutL3_43[2],gpcOutL3_114[1],gpcOutL3_115[0],gpcOutL3_136[2]},gpcOutL4_36);
wire [2:0] gpcOutL4_37;

// (* RLOC = "X4Y37" *)
gpc006 gpcL4_37 ({gpcOutL3_31[2],gpcOutL3_32[1],gpcOutL3_44[0],gpcOutL3_114[2],gpcOutL3_115[1],gpcOutL3_137[0]},gpcOutL4_37);
wire [2:0] gpcOutL4_38;

// (* RLOC = "X4Y38" *)
gpc006 gpcL4_38 ({gpcOutL3_32[2],gpcOutL3_33[0],gpcOutL3_44[1],gpcOutL3_115[2],gpcOutL3_116[0],gpcOutL3_137[1]},gpcOutL4_38);
wire [2:0] gpcOutL4_39;

// (* RLOC = "X4Y39" *)
gpc006 gpcL4_39 ({gpcOutL3_33[1],gpcOutL3_34[0],gpcOutL3_44[2],gpcOutL3_116[1],gpcOutL3_117[0],gpcOutL3_137[2]},gpcOutL4_39);
wire [2:0] gpcOutL4_40;

// (* RLOC = "X4Y40" *)
gpc006 gpcL4_40 ({gpcOutL3_24[2],gpcOutL3_25[1],gpcOutL3_35[0],gpcOutL3_93[2],gpcOutL3_94[1],gpcOutL3_118[0]},gpcOutL4_40);
wire [2:0] gpcOutL4_41;

// (* RLOC = "X4Y41" *)
gpc006 gpcL4_41 ({gpcOutL3_25[2],gpcOutL3_35[1],gpcOutL3_36[0],gpcOutL3_94[2],gpcOutL3_118[1],gpcOutL3_119[0]},gpcOutL4_41);
wire [2:0] gpcOutL4_42;

// (* RLOC = "X4Y42" *)
gpc006 gpcL4_42 ({gpcOutL3_35[2],gpcOutL3_36[1],gpcOutL3_37[0],gpcOutL3_118[2],gpcOutL3_119[1],gpcOutL3_120[0]},gpcOutL4_42);
wire [2:0] gpcOutL4_43;

// (* RLOC = "X4Y43" *)
gpc006 gpcL4_43 ({gpcOutL3_36[2],gpcOutL3_37[1],gpcOutL3_38[0],gpcOutL3_119[2],gpcOutL3_120[1],gpcOutL3_121[0]},gpcOutL4_43);
wire [2:0] gpcOutL4_44;

// (* RLOC = "X4Y44" *)
gpc006 gpcL4_44 ({gpcOutL3_37[2],gpcOutL3_38[1],gpcOutL3_39[0],gpcOutL3_120[2],gpcOutL3_121[1],gpcOutL3_122[0]},gpcOutL4_44);
wire [2:0] gpcOutL4_45;

// (* RLOC = "X4Y45" *)
gpc006 gpcL4_45 ({gpcOutL3_38[2],gpcOutL3_39[1],gpcOutL3_40[0],gpcOutL3_121[2],gpcOutL3_122[1],gpcOutL3_123[0]},gpcOutL4_45);
wire [2:0] gpcOutL4_46;

// (* RLOC = "X4Y46" *)
gpc006 gpcL4_46 ({gpcOutL3_30[1],gpcOutL3_40[2],gpcOutL3_46[0],gpcOutL3_108[1],gpcOutL3_123[2],gpcOutL3_139[0]},gpcOutL4_46);
wire [2:0] gpcOutL4_47;

// (* RLOC = "X4Y47" *)
gpc006 gpcL4_47 ({gpcOutL3_46[2],gpcOutL3_47[1],gpcOutL3_48[0],gpcOutL3_139[2],gpcOutL3_140[0],gpcOutL3_151[1]},gpcOutL4_47);
wire [2:0] gpcOutL4_48;

// (* RLOC = "X4Y48" *)
gpc006 gpcL4_48 ({gpcOutL3_47[2],gpcOutL3_48[1],gpcOutL3_49[0],gpcOutL3_140[1],gpcOutL3_152[0],pp63[26]},gpcOutL4_48);
wire [2:0] gpcOutL4_49;

// (* RLOC = "X4Y49" *)
gpc006 gpcL4_49 ({gpcOutL3_48[2],gpcOutL3_49[1],gpcOutL3_50[0],gpcOutL3_140[2],gpcOutL3_141[0],gpcOutL3_152[1]},gpcOutL4_49);
wire [2:0] gpcOutL4_50;

// (* RLOC = "X4Y50" *)
gpc006 gpcL4_50 ({gpcOutL3_49[2],gpcOutL3_50[1],gpcOutL3_76[0],gpcOutL3_141[1],gpcOutL2_272[1],gpcOutL2_290[0]},gpcOutL4_50);
wire [2:0] gpcOutL4_51;

// (* RLOC = "X4Y51" *)
gpc006 gpcL4_51 ({gpcOutL3_97[2],gpcOutL3_98[1],gpcOutL3_99[0],gpcOutL3_183[3],gpcOutL2_345[2],pp63[39]},gpcOutL4_51);
wire [2:0] gpcOutL4_52;

// (* RLOC = "X4Y52" *)
gpc015 gpcL4_52 ({gpcOutL3_82[1],gpcOutL3_82[0],gpcOutL3_112[2],gpcOutL3_113[1],pp24[1],pp25[0]},gpcOutL4_52);
wire [2:0] gpcOutL4_53;

// (* RLOC = "X4Y53" *)
gpc015 gpcL4_53 ({gpcOutL3_63[1],gpcOutL3_63[0],gpcOutL3_84[1],gpcOutL3_103[2],gpcOutL3_162[0],gpcOutL3_180[3]},gpcOutL4_53);
wire [2:0] gpcOutL4_54;

// (* RLOC = "X4Y54" *)
gpc015 gpcL4_54 ({gpcOutL3_41[0],gpcOutL3_65[1],gpcOutL3_66[0],gpcOutL3_85[2],gpcOutL3_163[1],gpcOutL2_320[1]},gpcOutL4_54);
wire [2:0] gpcOutL4_55;

// (* RLOC = "X4Y55" *)
gpc005 gpcL4_55 ({gpcOutL3_41[1],gpcOutL3_51[0],gpcOutL3_66[2],gpcOutL3_134[1],gpcOutL3_164[0]},gpcOutL4_55);
wire [2:0] gpcOutL4_56;

// (* RLOC = "X4Y56" *)
gpc005 gpcL4_56 ({gpcOutL3_51[2],gpcOutL3_52[1],gpcOutL3_53[0],gpcOutL3_146[1],gpcOutL3_165[0]},gpcOutL4_56);
wire [2:0] gpcOutL4_57;

// (* RLOC = "X4Y57" *)
gpc005 gpcL4_57 ({gpcOutL3_42[1],gpcOutL3_53[2],gpcOutL3_54[0],gpcOutL3_135[1],gpcOutL3_166[0]},gpcOutL4_57);
wire [2:0] gpcOutL4_58;

// (* RLOC = "X4Y58" *)
gpc005 gpcL4_58 ({gpcOutL3_31[0],gpcOutL3_43[1],gpcOutL3_54[2],gpcOutL3_114[0],gpcOutL3_136[1]},gpcOutL4_58);
wire [2:0] gpcOutL4_59;

// (* RLOC = "X4Y59" *)
gpc015 gpcL4_59 ({gpcOutL3_76[2],gpcOutL3_50[2],gpcOutL3_76[1],gpcOutL3_77[0],gpcOutL3_141[2],gpcOutL3_173[0]},gpcOutL4_59);
wire [2:0] gpcOutL4_60;

// (* RLOC = "X4Y60" *)
gpc015 gpcL4_60 ({gpcOutL3_78[2],gpcOutL3_77[2],gpcOutL3_78[1],gpcOutL3_79[0],gpcOutL3_173[2],gpcOutL3_174[0]},gpcOutL4_60);
wire [2:0] gpcOutL4_61;

// (* RLOC = "X4Y61" *)
gpc015 gpcL4_61 ({gpcOutL3_62[0],gpcOutL3_79[2],gpcOutL3_80[1],gpcOutL3_81[0],gpcOutL3_174[2],gpcOutL3_175[0]},gpcOutL4_61);
wire [2:0] gpcOutL4_62;

// (* RLOC = "X4Y62" *)
gpc015 gpcL4_62 ({gpcOutL3_62[2],gpcOutL3_62[1],gpcOutL3_81[2],gpcOutL3_95[0],gpcOutL3_153[1],gpcOutL2_344[0]},gpcOutL4_62);
wire [2:0] gpcOutL4_63;

// (* RLOC = "X4Y63" *)
gpc014 gpcL4_63 ({gpcOutL3_100[2],gpcOutL3_82[2],gpcOutL3_100[1],gpcOutL3_101[0],gpcOutL2_334[0]},gpcOutL4_63);
wire [2:0] gpcOutL4_64;

// (* RLOC = "X4Y64" *)
gpc014 gpcL4_64 ({gpcOutL3_83[1],gpcOutL3_83[0],gpcOutL3_101[2],gpcOutL3_102[1],gpcOutL3_180[0]},gpcOutL4_64);
wire [2:0] gpcOutL4_65;

// (* RLOC = "X4Y65" *)
gpc023 gpcL4_65 ({gpcOutL3_83[2],gpcOutL3_84[0],gpcOutL3_102[2],gpcOutL3_103[0],gpcOutL3_180[1]},gpcOutL4_65);
wire [1:0] gpcOutL4_66;

// (* RLOC = "X4Y66" *)
gpc003 gpcL4_66 ({gpcOutL3_64[0],gpcOutL3_84[2],gpcOutL3_162[1]},gpcOutL4_66);
wire [1:0] gpcOutL4_67;

// (* RLOC = "X4Y67" *)
gpc003 gpcL4_67 ({gpcOutL3_64[2],gpcOutL3_65[0],gpcOutL3_85[1]},gpcOutL4_67);
wire [1:0] gpcOutL4_68;

// (* RLOC = "X4Y68" *)
gpc003 gpcL4_68 ({gpcOutL3_65[2],gpcOutL3_66[1],gpcOutL3_134[0]},gpcOutL4_68);
wire [2:0] gpcOutL4_69;

// (* RLOC = "X4Y69" *)
gpc014 gpcL4_69 ({gpcOutL3_138[0],gpcOutL3_147[2],gpcOutL3_148[1],gpcOutL2_270[1],gpcOutL2_350[2]},gpcOutL4_69);
wire [1:0] gpcOutL4_70;

// (* RLOC = "X4Y70" *)
gpc003 gpcL4_70 ({gpcOutL3_77[1],gpcOutL3_78[0],gpcOutL3_173[1]},gpcOutL4_70);
wire [1:0] gpcOutL4_71;

// (* RLOC = "X4Y71" *)
gpc003 gpcL4_71 ({gpcOutL3_79[1],gpcOutL3_80[0],gpcOutL3_174[1]},gpcOutL4_71);
wire [1:0] gpcOutL4_72;

// (* RLOC = "X4Y72" *)
gpc003 gpcL4_72 ({gpcOutL3_80[2],gpcOutL3_81[1],gpcOutL3_153[0]},gpcOutL4_72);
wire [2:0] gpcOutL4_73;

// (* RLOC = "X4Y73" *)
gpc014 gpcL4_73 ({gpcOutL3_95[2],gpcOutL3_95[1],gpcOutL3_96[0],gpcOutL3_153[2],gpcOutL3_183[0]},gpcOutL4_73);
wire [2:0] gpcOutL4_74;

// (* RLOC = "X4Y74" *)
gpc023 gpcL4_74 ({gpcOutL3_96[2],gpcOutL3_97[1],gpcOutL3_96[1],gpcOutL3_97[0],gpcOutL3_183[1]},gpcOutL4_74);
wire [2:0] gpcOutL4_75;

// (* RLOC = "X4Y75" *)
gpc014 gpcL4_75 ({gpcOutL3_109[1],gpcOutL3_109[0],gpcOutL3_128[2],gpcOutL3_129[1],gpcOutL1_627[0]},gpcOutL4_75);
wire [2:0] gpcOutL4_76;

// (* RLOC = "X4Y76" *)
gpc014 gpcL4_76 ({gpcOutL3_142[2],gpcOutL3_109[2],gpcOutL3_142[1],gpcOutL3_154[0],gpcOutL1_669[0]},gpcOutL4_76);
wire [3:0] gpcOutL4_77;

// (* RLOC = "X4Y77" *)
gpc213 gpcL4_77 ({gpcOutL3_158[1],gpcOutL2_316[1],gpcOutL3_158[0],gpcOutL3_157[2],gpcOutL2_275[1],gpcOutL2_306[0]},gpcOutL4_77);
wire [2:0] gpcOutL4_78;

// (* RLOC = "X4Y78" *)
gpc023 gpcL4_78 ({gpcOutL3_145[1],gpcOutL3_160[0],gpcOutL3_130[2],gpcOutL3_145[0],gpcOutL3_159[1]},gpcOutL4_78);
wire [2:0] gpcOutL4_79;

// (* RLOC = "X4Y79" *)
gpc023 gpcL4_79 ({gpcOutL3_131[1],gpcOutL3_161[0],gpcOutL3_131[0],gpcOutL3_145[2],gpcOutL3_160[1]},gpcOutL4_79);
wire [2:0] gpcOutL4_80;

// (* RLOC = "X4Y80" *)
gpc023 gpcL4_80 ({gpcOutL3_110[0],gpcOutL3_132[1],gpcOutL3_131[2],gpcOutL3_132[0],gpcOutL3_161[1]},gpcOutL4_80);
wire [2:0] gpcOutL4_81;

// (* RLOC = "X4Y81" *)
gpc023 gpcL4_81 ({gpcOutL3_110[2],gpcOutL3_111[1],gpcOutL3_110[1],gpcOutL3_111[0],gpcOutL3_132[2]},gpcOutL4_81);
wire [2:0] gpcOutL4_82;

// (* RLOC = "X4Y82" *)
gpc023 gpcL4_82 ({gpcOutL3_112[1],gpcOutL3_113[0],gpcOutL3_111[2],gpcOutL3_112[0],gpcOutL3_133[1]},gpcOutL4_82);
wire [1:0] gpcOutL4_83;

// (* RLOC = "X4Y83" *)
gpc003 gpcL4_83 ({gpcOutL3_100[0],gpcOutL3_113[2],gpcOutL1_654[0]},gpcOutL4_83);
wire [1:0] gpcOutL4_84;

// (* RLOC = "X4Y84" *)
gpc003 gpcL4_84 ({gpcOutL3_101[1],gpcOutL3_102[0],gpcOutL2_334[1]},gpcOutL4_84);
wire [3:0] gpcOutL4_85;

// (* RLOC = "X4Y85" *)
gpc213 gpcL4_85 ({gpcOutL3_168[1],gpcOutL2_324[1],gpcOutL3_168[0],gpcOutL3_167[2],gpcOutL2_279[1],gpcOutL2_314[0]},gpcOutL4_85);
wire [2:0] gpcOutL4_86;

// (* RLOC = "X4Y86" *)
gpc023 gpcL4_86 ({gpcOutL3_149[1],gpcOutL3_170[0],gpcOutL3_138[2],gpcOutL3_149[0],gpcOutL3_169[1]},gpcOutL4_86);
wire [2:0] gpcOutL4_87;

// (* RLOC = "X4Y87" *)
gpc023 gpcL4_87 ({gpcOutL3_170[2],gpcOutL3_171[0],gpcOutL3_149[2],gpcOutL3_170[1],gpcOutL2_281[0]},gpcOutL4_87);
wire [1:0] gpcOutL4_88;

// (* RLOC = "X4Y88" *)
gpc003 gpcL4_88 ({gpcOutL3_182[3],gpcOutL2_341[2],pp63[15]},gpcOutL4_88);
wire [2:0] gpcOutL4_89;

// (* RLOC = "X4Y89" *)
gpc023 gpcL4_89 ({gpcOutL3_99[2],gpcOutL3_124[1],gpcOutL3_98[2],gpcOutL3_99[1],gpcOutL3_124[0]},gpcOutL4_89);
wire [2:0] gpcOutL4_90;

// (* RLOC = "X4Y90" *)
gpc023 gpcL4_90 ({gpcOutL3_125[2],gpcOutL3_126[1],gpcOutL3_124[2],gpcOutL3_125[1],gpcOutL3_126[0]},gpcOutL4_90);
wire [2:0] gpcOutL4_91;

// (* RLOC = "X4Y91" *)
gpc023 gpcL4_91 ({gpcOutL3_127[2],gpcOutL3_128[1],gpcOutL3_126[2],gpcOutL3_127[1],gpcOutL3_128[0]},gpcOutL4_91);
wire [2:0] gpcOutL4_92;

// (* RLOC = "X4Y92" *)
gpc023 gpcL4_92 ({gpcOutL3_143[2],gpcOutL3_144[0],gpcOutL3_143[1],gpcOutL3_155[0],pp63[50]},gpcOutL4_92);
wire [2:0] gpcOutL4_93;

// (* RLOC = "X4Y93" *)
gpc023 gpcL4_93 ({gpcOutL3_144[2],gpcOutL3_176[0],gpcOutL3_144[1],gpcOutL2_274[1],gpcOutL2_300[0]},gpcOutL4_93);
wire [1:0] gpcOutL4_94;

// (* RLOC = "X4Y94" *)
gpc003 gpcL4_94 ({gpcOutL3_184[3],gpcOutL2_349[2],pp63[63]},gpcOutL4_94);
wire [2:0] gpcOutL4_95;

// (* RLOC = "X4Y95" *)
gpc022 gpcL4_95 ({gpcOutL3_157[1],gpcOutL2_331[1],gpcOutL3_157[0],gpcOutL3_179[3]},gpcOutL4_95);
wire [2:0] gpcOutL4_96;

// (* RLOC = "X4Y96" *)
gpc022 gpcL4_96 ({gpcOutL3_130[1],gpcOutL3_159[0],gpcOutL3_130[0],gpcOutL3_158[2]},gpcOutL4_96);
wire [2:0] gpcOutL4_97;

// (* RLOC = "X4Y97" *)
gpc022 gpcL4_97 ({gpcOutL3_167[1],gpcOutL2_339[1],gpcOutL3_167[0],gpcOutL3_181[3]},gpcOutL4_97);
wire [2:0] gpcOutL4_98;

// (* RLOC = "X4Y98" *)
gpc022 gpcL4_98 ({gpcOutL3_147[1],gpcOutL3_148[0],gpcOutL3_147[0],gpcOutL3_168[2]},gpcOutL4_98);
wire [3:0] gpcOutL4_99;

// (* RLOC = "X4Y99" *)
gpc222 gpcL4_99 ({gpcOutL3_172[1],gpcOutL2_325[0],gpcOutL3_171[2],gpcOutL3_172[0],gpcOutL3_171[1],gpcOutL2_283[0]},gpcOutL4_99);
wire [3:0] gpcOutL4_100;

// (* RLOC = "X4Y100" *)
gpc222 gpcL4_100 ({gpcOutL3_150[2],gpcOutL3_182[0],gpcOutL3_150[1],gpcOutL2_340[0],gpcOutL3_150[0],gpcOutL3_172[2]},gpcOutL4_100);
wire [3:0] gpcOutL4_101;

// (* RLOC = "X4Y101" *)
gpc222 gpcL4_101 ({gpcOutL3_177[1],gpcOutL2_304[0],gpcOutL3_176[2],gpcOutL3_177[0],gpcOutL3_176[1],gpcOutL2_302[0]},gpcOutL4_101);
wire [3:0] gpcOutL4_102;

// (* RLOC = "X4Y102" *)
gpc222 gpcL4_102 ({gpcOutL3_156[1],gpcOutL2_348[0],gpcOutL3_156[0],gpcOutL3_178[1],gpcOutL3_177[2],gpcOutL3_178[0]},gpcOutL4_102);
wire [2:0] gpcOutL5_0;

// (* RLOC = "X5Y0" *)
gpc006 gpcL5_0 ({gpcOutL4_0[2],gpcOutL4_11[1],gpcOutL4_12[0],gpcOutL4_69[2],gpcOutL3_138[1],gpcOutL3_169[0]},gpcOutL5_0);
wire [2:0] gpcOutL5_1;

// (* RLOC = "X5Y1" *)
gpc015 gpcL5_1 ({gpcOutL4_5[1],gpcOutL4_5[0],gpcOutL4_38[2],gpcOutL4_39[1],pp48[1],pp49[0]},gpcOutL5_1);
wire [2:0] gpcOutL5_2;

// (* RLOC = "X5Y2" *)
gpc015 gpcL5_2 ({gpcOutL4_1[1],gpcOutL4_1[0],gpcOutL4_6[2],gpcOutL4_7[1],gpcOutL4_85[0],gpcOutL4_97[2]},gpcOutL5_2);
wire [2:0] gpcOutL5_3;

// (* RLOC = "X5Y3" *)
gpc015 gpcL5_3 ({gpcOutL4_8[2],gpcOutL4_8[1],gpcOutL4_9[0],gpcOutL4_27[2],gpcOutL4_85[3],gpcOutL4_98[0]},gpcOutL5_3);
wire [2:0] gpcOutL5_4;

// (* RLOC = "X5Y4" *)
gpc015 gpcL5_4 ({gpcOutL4_0[1],gpcOutL4_0[0],gpcOutL4_9[2],gpcOutL4_10[1],gpcOutL4_69[0],gpcOutL4_98[2]},gpcOutL5_4);
wire [2:0] gpcOutL5_5;

// (* RLOC = "X5Y5" *)
gpc015 gpcL5_5 ({gpcOutL4_3[1],gpcOutL4_2[2],gpcOutL4_3[0],gpcOutL4_13[1],gpcOutL4_86[2],gpcOutL4_87[0]},gpcOutL5_5);
wire [2:0] gpcOutL5_6;

// (* RLOC = "X5Y6" *)
gpc015 gpcL5_6 ({gpcOutL4_14[2],gpcOutL4_3[2],gpcOutL4_14[1],gpcOutL4_15[0],gpcOutL4_87[2],gpcOutL4_99[0]},gpcOutL5_6);
wire [2:0] gpcOutL5_7;

// (* RLOC = "X5Y7" *)
gpc015 gpcL5_7 ({gpcOutL4_17[2],gpcOutL4_16[2],gpcOutL4_17[1],gpcOutL4_18[0],gpcOutL4_99[3],gpcOutL4_100[0]},gpcOutL5_7);
wire [2:0] gpcOutL5_8;

// (* RLOC = "X5Y8" *)
gpc015 gpcL5_8 ({gpcOutL4_20[2],gpcOutL4_19[2],gpcOutL4_20[1],gpcOutL4_28[0],gpcOutL4_100[3],gpcOutL3_182[1]},gpcOutL5_8);
wire [2:0] gpcOutL5_9;

// (* RLOC = "X5Y9" *)
gpc014 gpcL5_9 ({gpcOutL4_53[0],gpcOutL4_64[2],gpcOutL4_65[1],gpcOutL3_103[1],gpcOutL3_180[2]},gpcOutL5_9);
wire [2:0] gpcOutL5_10;

// (* RLOC = "X5Y10" *)
gpc014 gpcL5_10 ({gpcOutL4_21[2],gpcOutL4_5[2],gpcOutL4_21[1],gpcOutL4_22[0],gpcOutL2_338[0]},gpcOutL5_10);
wire [2:0] gpcOutL5_11;

// (* RLOC = "X5Y11" *)
gpc014 gpcL5_11 ({gpcOutL4_23[2],gpcOutL4_22[2],gpcOutL4_23[1],gpcOutL4_24[0],gpcOutL3_181[0]},gpcOutL5_11);
wire [2:0] gpcOutL5_12;

// (* RLOC = "X5Y12" *)
gpc014 gpcL5_12 ({gpcOutL4_6[0],gpcOutL4_24[2],gpcOutL4_25[1],gpcOutL4_26[0],gpcOutL3_181[2]},gpcOutL5_12);
wire [2:0] gpcOutL5_13;

// (* RLOC = "X5Y13" *)
gpc023 gpcL5_13 ({gpcOutL4_6[1],gpcOutL4_7[0],gpcOutL4_25[2],gpcOutL4_26[1],gpcOutL4_97[0]},gpcOutL5_13);
wire [2:0] gpcOutL5_14;

// (* RLOC = "X5Y14" *)
gpc023 gpcL5_14 ({gpcOutL4_1[2],gpcOutL4_8[0],gpcOutL4_7[2],gpcOutL4_27[0],gpcOutL4_85[1]},gpcOutL5_14);
wire [1:0] gpcOutL5_15;

// (* RLOC = "X5Y15" *)
gpc003 gpcL5_15 ({gpcOutL4_10[2],gpcOutL4_11[0],gpcOutL4_69[1]},gpcOutL5_15);
wire [2:0] gpcOutL5_16;

// (* RLOC = "X5Y16" *)
gpc014 gpcL5_16 ({gpcOutL4_2[1],gpcOutL4_2[0],gpcOutL4_11[2],gpcOutL4_12[1],gpcOutL4_86[0]},gpcOutL5_16);
wire [2:0] gpcOutL5_17;

// (* RLOC = "X5Y17" *)
gpc023 gpcL5_17 ({gpcOutL4_15[2],gpcOutL4_16[1],gpcOutL4_15[1],gpcOutL4_16[0],gpcOutL4_99[1]},gpcOutL5_17);
wire [2:0] gpcOutL5_18;

// (* RLOC = "X5Y18" *)
gpc023 gpcL5_18 ({gpcOutL4_18[2],gpcOutL4_19[1],gpcOutL4_18[1],gpcOutL4_19[0],gpcOutL4_100[1]},gpcOutL5_18);
wire [2:0] gpcOutL5_19;

// (* RLOC = "X5Y19" *)
gpc014 gpcL5_19 ({gpcOutL4_4[1],gpcOutL4_4[0],gpcOutL4_28[2],gpcOutL4_29[1],gpcOutL4_88[0]},gpcOutL5_19);
wire [2:0] gpcOutL5_20;

// (* RLOC = "X5Y20" *)
gpc014 gpcL5_20 ({gpcOutL4_30[1],gpcOutL4_30[0],gpcOutL4_44[2],gpcOutL4_45[1],gpcOutL1_623[0]},gpcOutL5_20);
wire [2:0] gpcOutL5_21;

// (* RLOC = "X5Y21" *)
gpc014 gpcL5_21 ({gpcOutL4_31[1],gpcOutL4_30[2],gpcOutL4_31[0],gpcOutL4_46[1],gpcOutL1_665[0]},gpcOutL5_21);
wire [2:0] gpcOutL5_22;

// (* RLOC = "X5Y22" *)
gpc014 gpcL5_22 ({gpcOutL4_59[2],gpcOutL4_50[2],gpcOutL4_59[1],gpcOutL4_70[0],gpcOutL2_292[0]},gpcOutL5_22);
wire [2:0] gpcOutL5_23;

// (* RLOC = "X5Y23" *)
gpc014 gpcL5_23 ({gpcOutL4_51[0],gpcOutL4_73[2],gpcOutL4_74[1],gpcOutL3_98[0],gpcOutL3_183[2]},gpcOutL5_23);
wire [2:0] gpcOutL5_24;

// (* RLOC = "X5Y24" *)
gpc023 gpcL5_24 ({gpcOutL4_63[1],gpcOutL4_84[0],gpcOutL4_52[2],gpcOutL4_63[0],gpcOutL4_83[1]},gpcOutL5_24);
wire [2:0] gpcOutL5_25;

// (* RLOC = "X5Y25" *)
gpc023 gpcL5_25 ({gpcOutL4_64[1],gpcOutL4_65[0],gpcOutL4_63[2],gpcOutL4_64[0],gpcOutL4_84[1]},gpcOutL5_25);
wire [2:0] gpcOutL5_26;

// (* RLOC = "X5Y26" *)
gpc023 gpcL5_26 ({gpcOutL4_32[0],gpcOutL4_53[2],gpcOutL4_53[1],gpcOutL4_66[0],gpcOutL2_335[1]},gpcOutL5_26);
wire [2:0] gpcOutL5_27;

// (* RLOC = "X5Y27" *)
gpc023 gpcL5_27 ({gpcOutL4_32[2],gpcOutL4_54[0],gpcOutL4_32[1],gpcOutL4_67[0],gpcOutL3_163[0]},gpcOutL5_27);
wire [2:0] gpcOutL5_28;

// (* RLOC = "X5Y28" *)
gpc023 gpcL5_28 ({gpcOutL4_54[2],gpcOutL4_55[0],gpcOutL4_54[1],gpcOutL4_68[0],gpcOutL3_163[2]},gpcOutL5_28);
wire [2:0] gpcOutL5_29;

// (* RLOC = "X5Y29" *)
gpc023 gpcL5_29 ({gpcOutL4_33[2],gpcOutL4_34[0],gpcOutL4_33[1],gpcOutL4_55[2],gpcOutL4_56[0]},gpcOutL5_29);
wire [2:0] gpcOutL5_30;

// (* RLOC = "X5Y30" *)
gpc023 gpcL5_30 ({gpcOutL4_34[2],gpcOutL4_35[0],gpcOutL4_34[1],gpcOutL4_56[2],gpcOutL4_57[0]},gpcOutL5_30);
wire [2:0] gpcOutL5_31;

// (* RLOC = "X5Y31" *)
gpc023 gpcL5_31 ({gpcOutL4_35[2],gpcOutL4_36[0],gpcOutL4_35[1],gpcOutL4_57[2],gpcOutL4_58[0]},gpcOutL5_31);
wire [2:0] gpcOutL5_32;

// (* RLOC = "X5Y32" *)
gpc023 gpcL5_32 ({gpcOutL4_36[2],gpcOutL4_37[1],gpcOutL4_36[1],gpcOutL4_37[0],gpcOutL4_58[2]},gpcOutL5_32);
wire [1:0] gpcOutL5_33;

// (* RLOC = "X5Y33" *)
gpc003 gpcL5_33 ({gpcOutL4_37[2],gpcOutL4_38[1],gpcOutL4_39[0]},gpcOutL5_33);
wire [1:0] gpcOutL5_34;

// (* RLOC = "X5Y34" *)
gpc003 gpcL5_34 ({gpcOutL4_21[0],gpcOutL4_39[2],gpcOutL1_658[0]},gpcOutL5_34);
wire [1:0] gpcOutL5_35;

// (* RLOC = "X5Y35" *)
gpc003 gpcL5_35 ({gpcOutL4_22[1],gpcOutL4_23[0],gpcOutL2_338[1]},gpcOutL5_35);
wire [1:0] gpcOutL5_36;

// (* RLOC = "X5Y36" *)
gpc003 gpcL5_36 ({gpcOutL4_24[1],gpcOutL4_25[0],gpcOutL3_181[1]},gpcOutL5_36);
wire [1:0] gpcOutL5_37;

// (* RLOC = "X5Y37" *)
gpc003 gpcL5_37 ({gpcOutL4_9[1],gpcOutL4_10[0],gpcOutL4_98[1]},gpcOutL5_37);
wire [1:0] gpcOutL5_38;

// (* RLOC = "X5Y38" *)
gpc003 gpcL5_38 ({gpcOutL4_12[2],gpcOutL4_13[0],gpcOutL4_86[1]},gpcOutL5_38);
wire [1:0] gpcOutL5_39;

// (* RLOC = "X5Y39" *)
gpc003 gpcL5_39 ({gpcOutL4_13[2],gpcOutL4_14[0],gpcOutL4_87[1]},gpcOutL5_39);
wire [1:0] gpcOutL5_40;

// (* RLOC = "X5Y40" *)
gpc003 gpcL5_40 ({gpcOutL4_28[1],gpcOutL4_29[0],gpcOutL3_182[2]},gpcOutL5_40);
wire [2:0] gpcOutL5_41;

// (* RLOC = "X5Y41" *)
gpc023 gpcL5_41 ({gpcOutL4_4[2],gpcOutL4_40[1],gpcOutL4_29[2],gpcOutL4_40[0],gpcOutL4_88[1]},gpcOutL5_41);
wire [2:0] gpcOutL5_42;

// (* RLOC = "X5Y42" *)
gpc023 gpcL5_42 ({gpcOutL4_41[2],gpcOutL4_42[1],gpcOutL4_40[2],gpcOutL4_41[1],gpcOutL4_42[0]},gpcOutL5_42);
wire [2:0] gpcOutL5_43;

// (* RLOC = "X5Y43" *)
gpc023 gpcL5_43 ({gpcOutL4_43[2],gpcOutL4_44[1],gpcOutL4_42[2],gpcOutL4_43[1],gpcOutL4_44[0]},gpcOutL5_43);
wire [2:0] gpcOutL5_44;

// (* RLOC = "X5Y44" *)
gpc023 gpcL5_44 ({gpcOutL4_47[2],gpcOutL4_48[1],gpcOutL4_31[2],gpcOutL4_47[1],gpcOutL4_48[0]},gpcOutL5_44);
wire [2:0] gpcOutL5_45;

// (* RLOC = "X5Y45" *)
gpc023 gpcL5_45 ({gpcOutL4_49[2],gpcOutL4_50[1],gpcOutL4_48[2],gpcOutL4_49[1],gpcOutL4_50[0]},gpcOutL5_45);
wire [2:0] gpcOutL5_46;

// (* RLOC = "X5Y46" *)
gpc023 gpcL5_46 ({gpcOutL4_60[2],gpcOutL4_61[0],gpcOutL4_60[1],gpcOutL4_71[0],gpcOutL2_294[0]},gpcOutL5_46);
wire [2:0] gpcOutL5_47;

// (* RLOC = "X5Y47" *)
gpc023 gpcL5_47 ({gpcOutL4_61[2],gpcOutL4_62[0],gpcOutL4_61[1],gpcOutL4_72[0],gpcOutL3_175[1]},gpcOutL5_47);
wire [1:0] gpcOutL5_48;

// (* RLOC = "X5Y48" *)
gpc003 gpcL5_48 ({gpcOutL4_62[2],gpcOutL4_73[1],gpcOutL4_74[0]},gpcOutL5_48);
wire [2:0] gpcOutL5_49;

// (* RLOC = "X5Y49" *)
gpc023 gpcL5_49 ({gpcOutL4_89[2],gpcOutL4_90[0],gpcOutL4_51[2],gpcOutL4_89[1],gpcOutL3_125[0]},gpcOutL5_49);
wire [2:0] gpcOutL5_50;

// (* RLOC = "X5Y50" *)
gpc023 gpcL5_50 ({gpcOutL4_75[2],gpcOutL4_76[0],gpcOutL4_75[1],gpcOutL3_129[2],gpcOutL3_142[0]},gpcOutL5_50);
wire [2:0] gpcOutL5_51;

// (* RLOC = "X5Y51" *)
gpc023 gpcL5_51 ({gpcOutL4_76[2],gpcOutL4_92[0],gpcOutL4_76[1],gpcOutL3_143[0],gpcOutL3_154[1]},gpcOutL5_51);
wire [1:0] gpcOutL5_52;

// (* RLOC = "X5Y52" *)
gpc003 gpcL5_52 ({gpcOutL4_102[3],gpcOutL3_156[2],gpcOutL3_184[0]},gpcOutL5_52);
wire [3:0] gpcOutL5_53;

// (* RLOC = "X5Y53" *)
gpc212 gpcL5_53 ({gpcOutL4_78[0],gpcOutL4_96[2],gpcOutL4_96[1],gpcOutL4_77[3],gpcOutL4_96[0]},gpcOutL5_53);
wire [3:0] gpcOutL5_54;

// (* RLOC = "X5Y54" *)
gpc212 gpcL5_54 ({gpcOutL4_79[2],gpcOutL4_80[0],gpcOutL4_79[1],gpcOutL4_78[2],gpcOutL4_79[0]},gpcOutL5_54);
wire [3:0] gpcOutL5_55;

// (* RLOC = "X5Y55" *)
gpc222 gpcL5_55 ({gpcOutL4_81[2],gpcOutL4_82[0],gpcOutL4_81[1],gpcOutL3_133[0],gpcOutL4_80[2],gpcOutL4_81[0]},gpcOutL5_55);
wire [3:0] gpcOutL5_56;

// (* RLOC = "X5Y56" *)
gpc222 gpcL5_56 ({gpcOutL4_52[1],gpcOutL4_83[0],gpcOutL4_52[0],gpcOutL4_82[2],gpcOutL4_82[1],gpcOutL3_133[2]},gpcOutL5_56);
wire [3:0] gpcOutL5_57;

// (* RLOC = "X5Y57" *)
gpc222 gpcL5_57 ({gpcOutL4_91[1],gpcOutL3_129[0],gpcOutL4_90[2],gpcOutL4_91[0],gpcOutL4_90[1],gpcOutL3_127[0]},gpcOutL5_57);
wire [2:0] gpcOutL5_58;

// (* RLOC = "X5Y58" *)
gpc022 gpcL5_58 ({gpcOutL4_92[2],gpcOutL4_93[0],gpcOutL4_92[1],gpcOutL3_155[1]},gpcOutL5_58);
wire [2:0] gpcOutL6_0;

// (* RLOC = "X6Y0" *)
gpc014 gpcL6_0 ({gpcOutL5_2[0],gpcOutL5_12[2],gpcOutL5_13[1],gpcOutL4_26[2],gpcOutL4_97[1]},gpcOutL6_0);
wire [2:0] gpcOutL6_1;

// (* RLOC = "X6Y1" *)
gpc014 gpcL6_1 ({gpcOutL5_3[0],gpcOutL5_2[2],gpcOutL5_14[1],gpcOutL4_27[1],gpcOutL4_85[2]},gpcOutL6_1);
wire [2:0] gpcOutL6_2;

// (* RLOC = "X6Y2" *)
gpc014 gpcL6_2 ({gpcOutL5_7[0],gpcOutL5_6[2],gpcOutL5_17[1],gpcOutL4_17[0],gpcOutL4_99[2]},gpcOutL6_2);
wire [2:0] gpcOutL6_3;

// (* RLOC = "X6Y3" *)
gpc014 gpcL6_3 ({gpcOutL5_8[0],gpcOutL5_7[2],gpcOutL5_18[1],gpcOutL4_20[0],gpcOutL4_100[2]},gpcOutL6_3);
wire [3:0] gpcOutL6_4;

// (* RLOC = "X6Y4" *)
gpc213 gpcL6_4 ({gpcOutL5_29[1],gpcOutL4_56[1],gpcOutL5_29[0],gpcOutL5_28[2],gpcOutL4_33[0],gpcOutL4_55[1]},gpcOutL6_4);
wire [2:0] gpcOutL6_5;

// (* RLOC = "X6Y5" *)
gpc023 gpcL6_5 ({gpcOutL5_10[1],gpcOutL5_35[0],gpcOutL5_1[2],gpcOutL5_10[0],gpcOutL5_34[1]},gpcOutL6_5);
wire [2:0] gpcOutL6_6;

// (* RLOC = "X6Y6" *)
gpc023 gpcL6_6 ({gpcOutL5_11[1],gpcOutL5_36[0],gpcOutL5_10[2],gpcOutL5_11[0],gpcOutL5_35[1]},gpcOutL6_6);
wire [2:0] gpcOutL6_7;

// (* RLOC = "X6Y7" *)
gpc023 gpcL6_7 ({gpcOutL5_12[1],gpcOutL5_13[0],gpcOutL5_11[2],gpcOutL5_12[0],gpcOutL5_36[1]},gpcOutL6_7);
wire [2:0] gpcOutL6_8;

// (* RLOC = "X6Y8" *)
gpc023 gpcL6_8 ({gpcOutL5_4[1],gpcOutL5_15[0],gpcOutL5_3[2],gpcOutL5_4[0],gpcOutL5_37[1]},gpcOutL6_8);
wire [2:0] gpcOutL6_9;

// (* RLOC = "X6Y9" *)
gpc023 gpcL6_9 ({gpcOutL5_0[1],gpcOutL5_16[0],gpcOutL5_0[0],gpcOutL5_4[2],gpcOutL5_15[1]},gpcOutL6_9);
wire [2:0] gpcOutL6_10;

// (* RLOC = "X6Y10" *)
gpc023 gpcL6_10 ({gpcOutL5_5[0],gpcOutL5_16[2],gpcOutL5_0[2],gpcOutL5_16[1],gpcOutL5_38[0]},gpcOutL6_10);
wire [2:0] gpcOutL6_11;

// (* RLOC = "X6Y11" *)
gpc023 gpcL6_11 ({gpcOutL5_6[1],gpcOutL5_17[0],gpcOutL5_5[2],gpcOutL5_6[0],gpcOutL5_39[1]},gpcOutL6_11);
wire [2:0] gpcOutL6_12;

// (* RLOC = "X6Y12" *)
gpc023 gpcL6_12 ({gpcOutL5_19[1],gpcOutL5_41[0],gpcOutL5_8[2],gpcOutL5_19[0],gpcOutL5_40[1]},gpcOutL6_12);
wire [2:0] gpcOutL6_13;

// (* RLOC = "X6Y13" *)
gpc023 gpcL6_13 ({gpcOutL5_41[2],gpcOutL5_42[0],gpcOutL5_19[2],gpcOutL5_41[1],gpcOutL4_41[0]},gpcOutL6_13);
wire [2:0] gpcOutL6_14;

// (* RLOC = "X6Y14" *)
gpc023 gpcL6_14 ({gpcOutL5_20[2],gpcOutL5_21[0],gpcOutL5_20[1],gpcOutL4_45[2],gpcOutL4_46[0]},gpcOutL6_14);
wire [2:0] gpcOutL6_15;

// (* RLOC = "X6Y15" *)
gpc023 gpcL6_15 ({gpcOutL5_21[2],gpcOutL5_44[0],gpcOutL5_21[1],gpcOutL4_46[2],gpcOutL4_47[0]},gpcOutL6_15);
wire [2:0] gpcOutL6_16;

// (* RLOC = "X6Y16" *)
gpc023 gpcL6_16 ({gpcOutL5_22[2],gpcOutL5_46[0],gpcOutL5_22[1],gpcOutL4_60[0],gpcOutL4_70[1]},gpcOutL6_16);
wire [3:0] gpcOutL6_17;

// (* RLOC = "X6Y17" *)
gpc213 gpcL6_17 ({gpcOutL5_23[0],gpcOutL5_48[1],gpcOutL5_48[0],gpcOutL5_47[2],gpcOutL4_62[1],gpcOutL4_73[0]},gpcOutL6_17);
wire [3:0] gpcOutL6_18;

// (* RLOC = "X6Y18" *)
gpc132 gpcL6_18 ({gpcOutL5_49[0],gpcOutL5_23[2],gpcOutL4_51[1],gpcOutL4_89[0],gpcOutL5_23[1],gpcOutL4_74[2]},gpcOutL6_18);
wire [1:0] gpcOutL6_19;

// (* RLOC = "X6Y19" *)
gpc003 gpcL6_19 ({gpcOutL5_57[3],gpcOutL4_75[0],gpcOutL4_91[2]},gpcOutL6_19);
wire [3:0] gpcOutL6_20;

// (* RLOC = "X6Y20" *)
gpc212 gpcL6_20 ({gpcOutL5_24[2],gpcOutL5_25[0],gpcOutL5_24[1],gpcOutL5_24[0],gpcOutL5_56[3]},gpcOutL6_20);
wire [3:0] gpcOutL6_21;

// (* RLOC = "X6Y21" *)
gpc222 gpcL6_21 ({gpcOutL5_9[2],gpcOutL5_26[0],gpcOutL5_9[1],gpcOutL4_65[2],gpcOutL5_9[0],gpcOutL5_25[2]},gpcOutL6_21);
wire [3:0] gpcOutL6_22;

// (* RLOC = "X6Y22" *)
gpc222 gpcL6_22 ({gpcOutL5_27[1],gpcOutL4_67[1],gpcOutL5_26[2],gpcOutL5_27[0],gpcOutL5_26[1],gpcOutL4_66[1]},gpcOutL6_22);
wire [2:0] gpcOutL6_23;

// (* RLOC = "X6Y23" *)
gpc022 gpcL6_23 ({gpcOutL5_28[1],gpcOutL4_68[1],gpcOutL5_27[2],gpcOutL5_28[0]},gpcOutL6_23);
wire [3:0] gpcOutL6_24;

// (* RLOC = "X6Y24" *)
gpc222 gpcL6_24 ({gpcOutL5_30[2],gpcOutL5_31[0],gpcOutL5_30[1],gpcOutL4_57[1],gpcOutL5_29[2],gpcOutL5_30[0]},gpcOutL6_24);
wire [3:0] gpcOutL6_25;

// (* RLOC = "X6Y25" *)
gpc222 gpcL6_25 ({gpcOutL5_32[1],gpcOutL4_38[0],gpcOutL5_31[2],gpcOutL5_32[0],gpcOutL5_31[1],gpcOutL4_58[1]},gpcOutL6_25);
wire [3:0] gpcOutL6_26;

// (* RLOC = "X6Y26" *)
gpc222 gpcL6_26 ({gpcOutL5_1[1],gpcOutL5_34[0],gpcOutL5_1[0],gpcOutL5_33[1],gpcOutL5_32[2],gpcOutL5_33[0]},gpcOutL6_26);
wire [3:0] gpcOutL6_27;

// (* RLOC = "X6Y27" *)
gpc222 gpcL6_27 ({gpcOutL5_43[1],gpcOutL4_45[0],gpcOutL5_42[2],gpcOutL5_43[0],gpcOutL5_42[1],gpcOutL4_43[0]},gpcOutL6_27);
wire [3:0] gpcOutL6_28;

// (* RLOC = "X6Y28" *)
gpc222 gpcL6_28 ({gpcOutL5_45[1],gpcOutL4_59[0],gpcOutL5_44[2],gpcOutL5_45[0],gpcOutL5_44[1],gpcOutL4_49[0]},gpcOutL6_28);
wire [3:0] gpcOutL6_29;

// (* RLOC = "X6Y29" *)
gpc222 gpcL6_29 ({gpcOutL5_47[1],gpcOutL4_72[1],gpcOutL5_46[2],gpcOutL5_47[0],gpcOutL5_46[1],gpcOutL4_71[1]},gpcOutL6_29);
wire [3:0] gpcOutL6_30;

// (* RLOC = "X6Y30" *)
gpc212 gpcL6_30 ({gpcOutL5_51[2],gpcOutL5_58[0],gpcOutL5_51[1],gpcOutL5_50[2],gpcOutL5_51[0]},gpcOutL6_30);
wire [2:0] gpcOutL6_31;

// (* RLOC = "X6Y31" *)
gpc022 gpcL6_31 ({gpcOutL4_93[2],gpcOutL4_101[0],gpcOutL5_58[2],gpcOutL4_93[1]},gpcOutL6_31);
wire [127:0] adderIn0;
wire [127:0] adderIn1;
wire [127:0] adderIn2;
wire [128:0] adderOut;

assign adderIn0 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,gpcOutL5_45[2],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,gpcOutL5_43[2],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,gpcOutL5_40[0],1'b0,1'b0,gpcOutL5_18[0],1'b0,1'b0,1'b0,1'b0,gpcOutL5_39[0],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,gpcOutL5_37[0],1'b0,1'b0,gpcOutL5_14[0],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
assign adderIn1 = {1'b0,1'b0,1'b0,gpcOutL3_184[1],1'b0,1'b0,1'b0,gpcOutL4_102[0],1'b0,gpcOutL4_101[1],1'b0,1'b0,gpcOutL5_58[1],1'b0,1'b0,1'b0,1'b0,gpcOutL5_50[0],1'b0,1'b0,1'b0,gpcOutL5_57[0],gpcOutL5_49[1],1'b0,1'b0,gpcOutL6_18[0],1'b0,1'b0,gpcOutL6_29[3],1'b0,1'b0,gpcOutL6_29[0],1'b0,1'b0,gpcOutL5_22[0],1'b0,1'b0,gpcOutL6_28[0],1'b0,gpcOutL6_15[0],1'b0,1'b0,gpcOutL5_20[0],1'b0,1'b0,gpcOutL6_27[0],1'b0,gpcOutL6_13[0],1'b0,1'b0,gpcOutL5_8[1],gpcOutL5_18[2],1'b0,gpcOutL5_7[1],gpcOutL5_17[2],gpcOutL6_11[2],1'b0,1'b0,gpcOutL5_5[1],gpcOutL5_38[1],gpcOutL6_10[0],1'b0,gpcOutL6_9[0],gpcOutL3_148[2],1'b0,gpcOutL5_3[1],gpcOutL5_14[2],1'b0,gpcOutL5_2[1],gpcOutL5_13[2],gpcOutL6_7[2],1'b0,gpcOutL6_7[0],1'b0,gpcOutL6_6[0],1'b0,gpcOutL6_26[3],1'b0,1'b0,gpcOutL6_26[0],1'b0,1'b0,gpcOutL6_25[0],1'b0,1'b0,gpcOutL6_24[0],1'b0,1'b0,gpcOutL6_23[2],1'b0,gpcOutL6_23[0],1'b0,1'b0,gpcOutL6_22[0],1'b0,1'b0,1'b0,gpcOutL5_25[1],1'b0,1'b0,1'b0,1'b0,1'b0,gpcOutL5_56[0],1'b0,1'b0,1'b0,gpcOutL4_80[1],1'b0,1'b0,1'b0,gpcOutL4_78[1],1'b0,1'b0,1'b0,1'b0,1'b0,gpcOutL4_95[2],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,pp1[0],1'b0};
assign adderIn2 = {gpcOutL4_94[1],gpcOutL4_94[0],gpcOutL3_184[2],gpcOutL5_52[1],gpcOutL5_52[0],gpcOutL4_102[2],gpcOutL4_102[1],gpcOutL4_101[3],gpcOutL4_101[2],gpcOutL6_31[2],gpcOutL6_31[1],gpcOutL6_31[0],gpcOutL6_30[3],gpcOutL6_30[2],gpcOutL6_30[1],gpcOutL6_30[0],gpcOutL5_50[1],gpcOutL6_19[1],gpcOutL6_19[0],gpcOutL5_57[2],gpcOutL5_57[1],gpcOutL5_49[2],gpcOutL6_18[3],gpcOutL6_18[2],gpcOutL6_18[1],gpcOutL6_17[3],gpcOutL6_17[2],gpcOutL6_17[1],gpcOutL6_17[0],gpcOutL6_29[2],gpcOutL6_29[1],gpcOutL6_16[2],gpcOutL6_16[1],gpcOutL6_16[0],gpcOutL6_28[3],gpcOutL6_28[2],gpcOutL6_28[1],gpcOutL6_15[2],gpcOutL6_15[1],gpcOutL6_14[2],gpcOutL6_14[1],gpcOutL6_14[0],gpcOutL6_27[3],gpcOutL6_27[2],gpcOutL6_27[1],gpcOutL6_13[2],gpcOutL6_13[1],gpcOutL6_12[2],gpcOutL6_12[1],gpcOutL6_12[0],gpcOutL6_3[2],gpcOutL6_3[1],gpcOutL6_3[0],gpcOutL6_2[2],gpcOutL6_2[1],gpcOutL6_2[0],gpcOutL6_11[1],gpcOutL6_11[0],gpcOutL6_10[2],gpcOutL6_10[1],gpcOutL6_9[2],gpcOutL6_9[1],gpcOutL6_8[2],gpcOutL6_8[1],gpcOutL6_8[0],gpcOutL6_1[2],gpcOutL6_1[1],gpcOutL6_1[0],gpcOutL6_0[2],gpcOutL6_0[1],gpcOutL6_0[0],gpcOutL6_7[1],gpcOutL6_6[2],gpcOutL6_6[1],gpcOutL6_5[2],gpcOutL6_5[1],gpcOutL6_5[0],gpcOutL6_26[2],gpcOutL6_26[1],gpcOutL6_25[3],gpcOutL6_25[2],gpcOutL6_25[1],gpcOutL6_24[3],gpcOutL6_24[2],gpcOutL6_24[1],gpcOutL6_4[3],gpcOutL6_4[2],gpcOutL6_4[1],gpcOutL6_4[0],gpcOutL6_23[1],gpcOutL6_22[3],gpcOutL6_22[2],gpcOutL6_22[1],gpcOutL6_21[3],gpcOutL6_21[2],gpcOutL6_21[1],gpcOutL6_21[0],gpcOutL6_20[3],gpcOutL6_20[2],gpcOutL6_20[1],gpcOutL6_20[0],gpcOutL5_56[2],gpcOutL5_56[1],gpcOutL5_55[3],gpcOutL5_55[2],gpcOutL5_55[1],gpcOutL5_55[0],gpcOutL5_54[3],gpcOutL5_54[2],gpcOutL5_54[1],gpcOutL5_54[0],gpcOutL5_53[3],gpcOutL5_53[2],gpcOutL5_53[1],gpcOutL5_53[0],gpcOutL4_77[2],gpcOutL4_77[1],gpcOutL4_77[0],gpcOutL4_95[1],gpcOutL4_95[0],gpcOutL3_179[2],gpcOutL3_179[1],gpcOutL3_179[0],gpcOutL2_330[1],gpcOutL2_330[0],gpcOutL1_650[0],pp0[1],pp0[0]};
assign adderOut = adderIn0+ adderIn1+ adderIn2;
assign mult_out = adderOut;

endmodule
